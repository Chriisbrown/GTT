library ieee;
  use ieee.std_logic_1164.all;
  use ieee.std_logic_misc.all;
  use ieee.numeric_std.all;

  use work.Constants.all;
  use work.Types.all;
  package Arrays0 is

    constant initPredict : ty := to_ty(0);
    constant feature : intArray2D(nTrees-1 downto 0)(nNodes-1 downto 0) := ((4, 1, 0, 0, 1, 2, 3, -2, -2, -2, -2, -2, -2, -2, -2),
                (4, 1, 0, 3, 19, 0, 0, -2, -2, -2, -2, -2, -2, -2, -2),
                (1, 0, 4, 4, 4, 3, 0, -2, -2, -2, -2, -2, -2, -2, -2),
                (1, 0, 4, 4, 4, 3, 0, -2, -2, -2, -2, -2, -2, -2, -2),
                (4, 1, 0, 16, 17, 2, 3, -2, -2, -2, -2, -2, -2, -2, -2),
                (0, 1, 4, 4, 16, 1, 3, -2, -2, -2, -2, -2, -2, -2, -2),
                (0, 4, 1, 17, 2, 3, 1, -2, -2, -2, -2, -2, -2, -2, -2),
                (0, 1, 4, 18, 4, 17, 0, -2, -2, -2, -2, -2, -2, -2, -2),
                (4, 16, 2, 17, 18, 3, 0, -2, -2, -2, -2, -2, -2, -2, -2),
                (3, 2, 4, 1, 17, 12, 4, -2, -2, -2, -2, -2, -2, -2, -2),
                (1, 0, 1, 2, 3, 18, 16, -2, -2, -2, -2, -2, -2, -2, -2),
                (0, 4, 4, 10, 2, 20, 2, -2, -2, -2, -2, -2, -2, -2, -2),
                (18, 4, 18, 18, 0, 3, 4, -2, -2, -2, -2, -2, -2, -2, -2),
                (1, 2, 16, 3, 12, 0, 7, -2, -2, -2, -2, -2, -2, -2, -2),
                (1, 2, 17, 3, 5, 4, 18, -2, -2, -2, -2, -2, -2, -2, -2),
                (7, 17, 6, 5, 12, 20, 13, -2, -2, -2, -2, -2, -2, -2, -2),
                (0, 18, 18, 18, 4, 18, 4, -2, -2, -2, -2, -2, -2, -2, -2),
                (0, 4, 17, 0, 2, 7, 14, -2, -2, -2, -2, -2, -2, -2, -2),
                (18, 18, 4, 4, 2, 18, 2, -2, -2, -2, -2, -2, -2, -2, -2),
                (1, 17, 16, 7, 13, -2, 3, -2, -2, -2, -2, -2, -2, -2, -2),
                (1, 5, 17, 8, 2, 7, 12, -2, -2, -2, -2, -2, -2, -2, -2),
                (3, 2, 1, 1, 17, 8, 16, -2, -2, -2, -2, -2, -2, -2, -2),
                (2, 3, 17, 18, 2, 6, 16, -2, -2, -2, -2, -2, -2, -2, -2),
                (0, 2, 1, 6, 17, 5, 16, -2, -2, -2, -2, -2, -2, -2, -2),
                (18, 4, 18, 3, -2, 3, 20, -2, -2, -2, -2, -2, -2, -2, -2),
                (1, 16, 17, 7, 4, 6, 19, -2, -2, -2, -2, -2, -2, -2, -2),
                (17, 7, 12, 5, 6, 17, 15, -2, -2, -2, -2, -2, -2, -2, -2),
                (2, 18, 17, 4, 18, -2, 3, -2, -2, -2, -2, -2, -2, -2, -2),
                (2, 17, 16, 6, 3, -2, 16, -2, -2, -2, -2, -2, -2, -2, -2),
                (0, -2, 3, 17, 3, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2),
                (18, 17, 16, 4, -2, 7, 4, -2, -2, -2, -2, -2, -2, -2, -2),
                (17, 7, 13, 5, 13, 5, 12, -2, -2, -2, -2, -2, -2, -2, -2),
                (0, 6, 17, 17, 17, 8, 16, -2, -2, -2, -2, -2, -2, -2, -2),
                (17, 5, 19, 9, 4, 10, 17, -2, -2, -2, -2, -2, -2, -2, -2),
                (18, 19, 18, 7, 5, 10, 4, -2, -2, -2, -2, -2, -2, -2, -2),
                (3, 2, 2, 16, 10, 3, 16, -2, -2, -2, -2, -2, -2, -2, -2),
                (1, 0, 16, -2, 3, 2, 7, -2, -2, -2, -2, -2, -2, -2, -2),
                (7, 13, 13, 10, 12, 6, 19, -2, -2, -2, -2, -2, -2, -2, -2),
                (16, 2, 16, 4, -2, 3, 4, -2, -2, -2, -2, -2, -2, -2, -2),
                (1, 16, 15, 2, 4, 17, 17, -2, -2, -2, -2, -2, -2, -2, -2),
                (7, 13, 13, 10, 12, 10, 4, -2, -2, -2, -2, -2, -2, -2, -2),
                (2, 1, 16, 16, 16, 16, 16, -2, -2, -2, -2, -2, -2, -2, -2),
                (18, 0, 3, 4, 18, 4, -2, -2, -2, -2, -2, -2, -2, -2, -2),
                (0, 17, 3, -2, 16, 1, 3, -2, -2, -2, -2, -2, -2, -2, -2),
                (0, 5, 16, 8, 16, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2),
                (17, 20, 14, 6, 2, 15, 19, -2, -2, -2, -2, -2, -2, -2, -2),
                (17, 8, 4, 16, 16, 16, 16, -2, -2, -2, -2, -2, -2, -2, -2),
                (18, 3, 16, 16, -2, 1, 4, -2, -2, -2, -2, -2, -2, -2, -2),
                (16, 2, 17, 4, -2, 7, 14, -2, -2, -2, -2, -2, -2, -2, -2),
                (18, 18, 4, 17, 5, 0, 16, -2, -2, -2, -2, -2, -2, -2, -2)
                );
    constant threshold_int : intArray2D(nTrees-1 downto 0)(nNodes-1 downto 0) := ((576, 2, 2112, 1856, 4, 8, 8, 0, 0, 0, 0, 0, 0, 0, 0),
                (576, 2, 1984, 6, 320, 1600, 2368, 0, 0, 0, 0, 0, 0, 0, 0),
                (4, 1856, 704, 576, 576, 4, 1984, 0, 0, 0, 0, 0, 0, 0, 0),
                (2, 1728, 704, 576, 704, 6, 1856, 0, 0, 0, 0, 0, 0, 0, 0),
                (576, 2, 1984, 18, 411, 8, 8, 0, 0, 0, 0, 0, 0, 0, 0),
                (1472, 4, 704, 576, 38, 2, 8, 0, 0, 0, 0, 0, 0, 0, 0),
                (1600, 576, 4, 116, 8, 6, 4, 0, 0, 0, 0, 0, 0, 0, 0),
                (1344, 4, 704, 40, 576, 396, 2240, 0, 0, 0, 0, 0, 0, 0, 0),
                (576, 26, 8, 134, -36, 8, 2240, 0, 0, 0, 0, 0, 0, 0, 0),
                (6, 6, 576, 4, 449, 64, 704, 0, 0, 0, 0, 0, 0, 0, 0),
                (2, 1216, 4, 4, 8, 39, 36, 0, 0, 0, 0, 0, 0, 0, 0),
                (1088, 576, 704, 64, 6, 192, 10, 0, 0, 0, 0, 0, 0, 0, 0),
                (-35, 576, 32, -42, 1600, 6, 576, 0, 0, 0, 0, 0, 0, 0, 0),
                (4, 10, 44, 8, 64, 448, 64, 0, 0, 0, 0, 0, 0, 0, 0),
                (2, 8, 109, 8, 64, 704, -28, 0, 0, 0, 0, 0, 0, 0, 0),
                (64, 294, 64, 64, 64, 576, 64, 0, 0, 0, 0, 0, 0, 0, 0),
                (960, 38, 44, -27, 576, -42, 704, 0, 0, 0, 0, 0, 0, 0, 0),
                (1088, 576, 557, 704, 6, 64, 64, 0, 0, 0, 0, 0, 0, 0, 0),
                (24, -23, 704, 576, 12, 44, 8, 0, 0, 0, 0, 0, 0, 0, 0),
                (4, 391, 36, 64, 64, 0, 4, 0, 0, 0, 0, 0, 0, -256, -256),
                (0, 64, 265, 64, 10, 64, 64, 0, 0, 0, 0, 0, 0, 0, 0),
                (6, 4, 2, 4, 262, 64, 22, 0, 0, 0, 0, 0, 0, 0, 0),
                (12, 8, 266, 38, 6, 64, 8, 0, 0, 0, 0, 0, 0, 0, 0),
                (832, 2, 4, 64, 78, 64, 34, 0, 0, 0, 0, 0, 0, 0, 0),
                (-42, 704, 24, 8, 0, 8, 576, 0, 0, 0, 0, 0, 0, -256, -256),
                (0, 28, 92, 64, 576, 64, 192, 0, 0, 0, 0, 0, 0, 0, 0),
                (283, 64, 64, 64, 64, 346, 64, 0, 0, 0, 0, 0, 0, 0, 0),
                (12, -29, 257, 576, 48, 0, 6, 0, 0, 0, 0, 0, 0, -256, -256),
                (12, 545, 2, 64, 6, 0, 32, 0, 0, 0, 0, 0, 0, -256, -256),
                (576, 0, 2, 247, 6, 0, 0, 0, 0, -256, -256, -256, -256, -256, -256),
                (-52, 519, 46, 704, 0, 64, 576, 0, 0, 0, 0, 0, 0, -256, -256),
                (376, 64, 64, 64, 64, 64, 64, 0, 0, 0, 0, 0, 0, 0, 0),
                (832, 64, 246, 551, 195, 64, 14, 0, 0, 0, 0, 0, 0, 0, 0),
                (72, 64, 192, 64, 704, 64, 269, 0, 0, 0, 0, 0, 0, 0, 0),
                (-18, 320, 20, 64, 64, 64, 576, 0, 0, 0, 0, 0, 0, 0, 0),
                (6, 8, 6, 6, 64, 8, 30, 0, 0, 0, 0, 0, 0, 0, 0),
                (4, 576, 34, 0, 4, 10, 64, 0, 0, 0, 0, 0, 0, -256, -256),
                (64, 64, 64, 64, 64, 64, 320, 0, 0, 0, 0, 0, 0, 0, 0),
                (0, 8, 46, 576, 0, 8, 576, 0, 0, 0, 0, 0, 0, -256, -256),
                (0, 24, 64, 10, 576, 376, 355, 0, 0, 0, 0, 0, 0, 0, 0),
                (64, 64, 64, 64, 64, 64, 576, 0, 0, 0, 0, 0, 0, 0, 0),
                (12, 4, 26, 38, 32, 10, 42, 0, 0, 0, 0, 0, 0, 0, 0),
                (52, 1088, 10, 704, -18, 704, 0, 0, 0, 0, 0, 0, 0, -256, -256),
                (704, 42, 2, 0, 30, 2, 6, 0, 0, 0, 0, 0, 0, -256, -256),
                (2624, 64, 42, 64, 30, 0, 0, 0, 0, 0, 0, -256, -256, -256, -256),
                (250, 320, 64, 64, 8, 64, 320, 0, 0, 0, 0, 0, 0, 0, 0),
                (60, 64, 576, 38, 24, 14, 32, 0, 0, 0, 0, 0, 0, 0, 0),
                (-52, 8, 46, 46, 0, 6, 576, 0, 0, 0, 0, 0, 0, -256, -256),
                (0, 8, 308, 576, 0, 64, 64, 0, 0, 0, 0, 0, 0, -256, -256),
                (20, -18, 576, 39, 64, 1856, 20, 0, 0, 0, 0, 0, 0, 0, 0)
                );
    constant children_left : intArray2D(nTrees-1 downto 0)(nNodes-1 downto 0) := ((1, 3, 5, 7, 9, 11, 13, -1, -1, -1, -1, -1, -1, -1, -1),
                (1, 3, 5, 7, 9, 11, 13, -1, -1, -1, -1, -1, -1, -1, -1),
                (1, 3, 5, 7, 9, 11, 13, -1, -1, -1, -1, -1, -1, -1, -1),
                (1, 3, 5, 7, 9, 11, 13, -1, -1, -1, -1, -1, -1, -1, -1),
                (1, 3, 5, 7, 9, 11, 13, -1, -1, -1, -1, -1, -1, -1, -1),
                (1, 3, 5, 7, 9, 11, 13, -1, -1, -1, -1, -1, -1, -1, -1),
                (1, 3, 5, 7, 9, 11, 13, -1, -1, -1, -1, -1, -1, -1, -1),
                (1, 3, 5, 7, 9, 11, 13, -1, -1, -1, -1, -1, -1, -1, -1),
                (1, 3, 5, 7, 9, 11, 13, -1, -1, -1, -1, -1, -1, -1, -1),
                (1, 3, 5, 7, 9, 11, 13, -1, -1, -1, -1, -1, -1, -1, -1),
                (1, 3, 5, 7, 9, 11, 13, -1, -1, -1, -1, -1, -1, -1, -1),
                (1, 3, 5, 7, 9, 11, 13, -1, -1, -1, -1, -1, -1, -1, -1),
                (1, 3, 5, 7, 9, 11, 13, -1, -1, -1, -1, -1, -1, -1, -1),
                (1, 3, 5, 7, 9, 11, 13, -1, -1, -1, -1, -1, -1, -1, -1),
                (1, 3, 5, 7, 9, 11, 13, -1, -1, -1, -1, -1, -1, -1, -1),
                (1, 3, 5, 7, 9, 11, 13, -1, -1, -1, -1, -1, -1, -1, -1),
                (1, 3, 5, 7, 9, 11, 13, -1, -1, -1, -1, -1, -1, -1, -1),
                (1, 3, 5, 7, 9, 11, 13, -1, -1, -1, -1, -1, -1, -1, -1),
                (1, 3, 5, 7, 9, 11, 13, -1, -1, -1, -1, -1, -1, -1, -1),
                (1, 3, 5, 7, 9, 13, 11, -1, -1, -1, -1, -1, -1, -1, -1),
                (1, 3, 5, 7, 9, 11, 13, -1, -1, -1, -1, -1, -1, -1, -1),
                (1, 3, 5, 7, 9, 11, 13, -1, -1, -1, -1, -1, -1, -1, -1),
                (1, 3, 5, 7, 9, 11, 13, -1, -1, -1, -1, -1, -1, -1, -1),
                (1, 3, 5, 7, 9, 11, 13, -1, -1, -1, -1, -1, -1, -1, -1),
                (1, 3, 5, 7, 13, 9, 11, -1, -1, -1, -1, -1, -1, -1, -1),
                (1, 3, 5, 7, 9, 11, 13, -1, -1, -1, -1, -1, -1, -1, -1),
                (1, 3, 5, 7, 9, 11, 13, -1, -1, -1, -1, -1, -1, -1, -1),
                (1, 3, 5, 7, 9, 13, 11, -1, -1, -1, -1, -1, -1, -1, -1),
                (1, 3, 5, 7, 9, 13, 11, -1, -1, -1, -1, -1, -1, -1, -1),
                (1, 9, 3, 5, 7, -1, -1, -1, -1, 11, 13, -1, -1, -1, -1),
                (1, 3, 5, 7, 13, 9, 11, -1, -1, -1, -1, -1, -1, -1, -1),
                (1, 3, 5, 7, 9, 11, 13, -1, -1, -1, -1, -1, -1, -1, -1),
                (1, 3, 5, 7, 9, 11, 13, -1, -1, -1, -1, -1, -1, -1, -1),
                (1, 3, 5, 7, 9, 11, 13, -1, -1, -1, -1, -1, -1, -1, -1),
                (1, 3, 5, 7, 9, 11, 13, -1, -1, -1, -1, -1, -1, -1, -1),
                (1, 3, 5, 7, 9, 11, 13, -1, -1, -1, -1, -1, -1, -1, -1),
                (1, 3, 5, 13, 7, 9, 11, -1, -1, -1, -1, -1, -1, -1, -1),
                (1, 3, 5, 7, 9, 11, 13, -1, -1, -1, -1, -1, -1, -1, -1),
                (1, 3, 5, 7, 13, 9, 11, -1, -1, -1, -1, -1, -1, -1, -1),
                (1, 3, 5, 7, 9, 11, 13, -1, -1, -1, -1, -1, -1, -1, -1),
                (1, 3, 5, 7, 9, 11, 13, -1, -1, -1, -1, -1, -1, -1, -1),
                (1, 3, 5, 7, 9, 11, 13, -1, -1, -1, -1, -1, -1, -1, -1),
                (1, 3, 5, 7, 9, 11, 13, -1, -1, -1, -1, -1, -1, -1, -1),
                (1, 3, 5, 13, 7, 9, 11, -1, -1, -1, -1, -1, -1, -1, -1),
                (1, 3, 5, 7, 9, 11, 13, -1, -1, -1, -1, -1, -1, -1, -1),
                (1, 3, 5, 7, 9, 11, 13, -1, -1, -1, -1, -1, -1, -1, -1),
                (1, 3, 5, 7, 9, 11, 13, -1, -1, -1, -1, -1, -1, -1, -1),
                (1, 3, 5, 7, 13, 9, 11, -1, -1, -1, -1, -1, -1, -1, -1),
                (1, 3, 5, 7, 13, 9, 11, -1, -1, -1, -1, -1, -1, -1, -1),
                (1, 3, 5, 7, 9, 11, 13, -1, -1, -1, -1, -1, -1, -1, -1)
                );
    constant children_right : intArray2D(nTrees-1 downto 0)(nNodes-1 downto 0) := ((2, 4, 6, 8, 10, 12, 14, -1, -1, -1, -1, -1, -1, -1, -1),
                (2, 4, 6, 8, 10, 12, 14, -1, -1, -1, -1, -1, -1, -1, -1),
                (2, 4, 6, 8, 10, 12, 14, -1, -1, -1, -1, -1, -1, -1, -1),
                (2, 4, 6, 8, 10, 12, 14, -1, -1, -1, -1, -1, -1, -1, -1),
                (2, 4, 6, 8, 10, 12, 14, -1, -1, -1, -1, -1, -1, -1, -1),
                (2, 4, 6, 8, 10, 12, 14, -1, -1, -1, -1, -1, -1, -1, -1),
                (2, 4, 6, 8, 10, 12, 14, -1, -1, -1, -1, -1, -1, -1, -1),
                (2, 4, 6, 8, 10, 12, 14, -1, -1, -1, -1, -1, -1, -1, -1),
                (2, 4, 6, 8, 10, 12, 14, -1, -1, -1, -1, -1, -1, -1, -1),
                (2, 4, 6, 8, 10, 12, 14, -1, -1, -1, -1, -1, -1, -1, -1),
                (2, 4, 6, 8, 10, 12, 14, -1, -1, -1, -1, -1, -1, -1, -1),
                (2, 4, 6, 8, 10, 12, 14, -1, -1, -1, -1, -1, -1, -1, -1),
                (2, 4, 6, 8, 10, 12, 14, -1, -1, -1, -1, -1, -1, -1, -1),
                (2, 4, 6, 8, 10, 12, 14, -1, -1, -1, -1, -1, -1, -1, -1),
                (2, 4, 6, 8, 10, 12, 14, -1, -1, -1, -1, -1, -1, -1, -1),
                (2, 4, 6, 8, 10, 12, 14, -1, -1, -1, -1, -1, -1, -1, -1),
                (2, 4, 6, 8, 10, 12, 14, -1, -1, -1, -1, -1, -1, -1, -1),
                (2, 4, 6, 8, 10, 12, 14, -1, -1, -1, -1, -1, -1, -1, -1),
                (2, 4, 6, 8, 10, 12, 14, -1, -1, -1, -1, -1, -1, -1, -1),
                (2, 4, 6, 8, 10, 14, 12, -1, -1, -1, -1, -1, -1, -1, -1),
                (2, 4, 6, 8, 10, 12, 14, -1, -1, -1, -1, -1, -1, -1, -1),
                (2, 4, 6, 8, 10, 12, 14, -1, -1, -1, -1, -1, -1, -1, -1),
                (2, 4, 6, 8, 10, 12, 14, -1, -1, -1, -1, -1, -1, -1, -1),
                (2, 4, 6, 8, 10, 12, 14, -1, -1, -1, -1, -1, -1, -1, -1),
                (2, 4, 6, 8, 14, 10, 12, -1, -1, -1, -1, -1, -1, -1, -1),
                (2, 4, 6, 8, 10, 12, 14, -1, -1, -1, -1, -1, -1, -1, -1),
                (2, 4, 6, 8, 10, 12, 14, -1, -1, -1, -1, -1, -1, -1, -1),
                (2, 4, 6, 8, 10, 14, 12, -1, -1, -1, -1, -1, -1, -1, -1),
                (2, 4, 6, 8, 10, 14, 12, -1, -1, -1, -1, -1, -1, -1, -1),
                (2, 10, 4, 6, 8, -1, -1, -1, -1, 12, 14, -1, -1, -1, -1),
                (2, 4, 6, 8, 14, 10, 12, -1, -1, -1, -1, -1, -1, -1, -1),
                (2, 4, 6, 8, 10, 12, 14, -1, -1, -1, -1, -1, -1, -1, -1),
                (2, 4, 6, 8, 10, 12, 14, -1, -1, -1, -1, -1, -1, -1, -1),
                (2, 4, 6, 8, 10, 12, 14, -1, -1, -1, -1, -1, -1, -1, -1),
                (2, 4, 6, 8, 10, 12, 14, -1, -1, -1, -1, -1, -1, -1, -1),
                (2, 4, 6, 8, 10, 12, 14, -1, -1, -1, -1, -1, -1, -1, -1),
                (2, 4, 6, 14, 8, 10, 12, -1, -1, -1, -1, -1, -1, -1, -1),
                (2, 4, 6, 8, 10, 12, 14, -1, -1, -1, -1, -1, -1, -1, -1),
                (2, 4, 6, 8, 14, 10, 12, -1, -1, -1, -1, -1, -1, -1, -1),
                (2, 4, 6, 8, 10, 12, 14, -1, -1, -1, -1, -1, -1, -1, -1),
                (2, 4, 6, 8, 10, 12, 14, -1, -1, -1, -1, -1, -1, -1, -1),
                (2, 4, 6, 8, 10, 12, 14, -1, -1, -1, -1, -1, -1, -1, -1),
                (2, 4, 6, 8, 10, 12, 14, -1, -1, -1, -1, -1, -1, -1, -1),
                (2, 4, 6, 14, 8, 10, 12, -1, -1, -1, -1, -1, -1, -1, -1),
                (2, 4, 6, 8, 10, 12, 14, -1, -1, -1, -1, -1, -1, -1, -1),
                (2, 4, 6, 8, 10, 12, 14, -1, -1, -1, -1, -1, -1, -1, -1),
                (2, 4, 6, 8, 10, 12, 14, -1, -1, -1, -1, -1, -1, -1, -1),
                (2, 4, 6, 8, 14, 10, 12, -1, -1, -1, -1, -1, -1, -1, -1),
                (2, 4, 6, 8, 14, 10, 12, -1, -1, -1, -1, -1, -1, -1, -1),
                (2, 4, 6, 8, 10, 12, 14, -1, -1, -1, -1, -1, -1, -1, -1)
                );
    constant value_int : intArray2D(nTrees-1 downto 0)(nNodes-1 downto 0) := ((0, 0, 0, 0, 0, 0, 0, 39, -24, -33, -62, 69, 50, 16, -35),
                (0, 0, 0, 0, 0, 0, 0, 27, -25, -46, -6, 54, 41, 17, -30),
                (0, 0, 0, 0, 0, 0, 0, 20, 45, -21, 17, -25, -45, 36, -15),
                (0, 0, 0, 0, 0, 0, 0, 23, 41, -3, 27, -12, -39, 37, 0),
                (0, 0, 0, 0, 0, 0, 0, -12, 25, -28, 14, 39, 24, 9, -24),
                (0, 0, 0, 0, 0, 0, 0, 21, 36, -33, 1, 6, -21, 25, -19),
                (0, 0, 0, 0, 0, 0, 0, -14, 20, 34, 18, 10, -15, -17, -37),
                (0, 0, 0, 0, 0, 0, 0, 30, -9, -14, 25, -14, 17, 21, -7),
                (0, 0, 0, 0, 0, 0, 0, -30, -11, -35, 11, 28, -28, 9, -10),
                (0, 0, 0, 0, 0, 0, 0, 27, -3, -1, 26, -29, -10, -11, 1),
                (0, 0, 0, 0, 0, 0, 0, 30, 18, 11, -10, 0, -34, -33, -5),
                (0, 0, 0, 0, 0, 0, 0, 19, -20, 29, 6, 13, -9, 19, 2),
                (0, 0, 0, 0, 0, 0, 0, -39, -22, 8, -13, 10, -8, -31, 0),
                (0, 0, 0, 0, 0, 0, 0, 10, -11, -15, 0, 0, -26, 0, 16),
                (0, 0, 0, 0, 0, 0, 0, 17, -17, 16, 0, -22, 10, -18, 2),
                (0, 0, 0, 0, 0, 0, 0, 14, -49, -28, 11, -28, 0, 14, -7),
                (0, 0, 0, 0, 0, 0, 0, 1, 21, -18, 0, -27, 1, -32, 0),
                (0, 0, 0, 0, 0, 0, 0, 19, -2, 21, 0, -10, 2, 29, 5),
                (0, 0, 0, 0, 0, 0, 0, -15, 0, 6, -6, -11, -28, 17, 0),
                (0, 0, 0, 0, 0, -23, 0, -15, 4, -23, 12, 7, -5, -23, -23),
                (0, 0, 0, 0, 0, 0, 0, 7, 33, 10, 2, -30, 0, -17, 7),
                (0, 0, 0, 0, 0, 0, 0, 17, 0, -3, 7, -6, 3, -18, -6),
                (0, 0, 0, 0, 0, 0, 0, 3, -15, -28, -5, 0, -22, -19, -3),
                (0, 0, 0, 0, 0, 0, 0, 0, 23, 0, 11, 6, -1, -19, 0),
                (0, 0, 0, 0, 0, 0, 0, -22, 0, 2, -10, -10, 6, 0, 0),
                (0, 0, 0, 0, 0, 0, 0, 2, 13, 8, -3, -27, -2, 5, -2),
                (0, 0, 0, 0, 0, 0, 0, 31, -31, -15, 3, 6, -23, 13, -1),
                (0, 0, 0, 0, 0, -18, 0, -13, 0, 2, -19, 0, -13, -18, -18),
                (0, 0, 0, 0, 0, -31, 0, -8, 1, 13, 0, -2, -16, -31, -31),
                (0, 18, 0, 0, 0, -13, 2, 2, -2, 18, 18, 18, 18, 18, 18),
                (0, 0, 0, 0, 0, 0, 0, -27, 0, -3, 1, 23, -7, 0, 0),
                (0, 0, 0, 0, 0, 0, 0, 13, -13, 3, -11, -36, -8, -15, 9),
                (0, 0, 0, 0, 0, 0, 0, -5, 9, 17, 0, -11, 1, -6, 4),
                (0, 0, 0, 0, 0, 0, 0, -20, 15, -15, 4, 9, -5, -8, 1),
                (0, 0, 0, 0, 0, 0, 0, -14, -3, -6, 3, 3, -1, -7, 1),
                (0, 0, 0, 0, 0, 0, 0, 25, 1, 1, -11, -4, -21, -5, 2),
                (0, 0, 0, 14, 0, 0, 0, -3, 1, -18, -6, -4, 5, 14, 14),
                (0, 0, 0, 0, 0, 0, 0, -18, 1, -9, 4, -8, 4, -22, 0),
                (0, 0, 0, 0, -41, 0, 0, 0, 23, 0, -7, 17, -8, -41, -41),
                (0, 0, 0, 0, 0, 0, 0, 11, 0, 6, -2, -1, 9, 19, -7),
                (0, 0, 0, 0, 0, 0, 0, -13, 0, -8, 3, 5, -2, -22, 0),
                (0, 0, 0, 0, 0, 0, 0, 2, -1, -11, 0, -10, 0, -22, 0),
                (0, 0, 0, 0, 0, 0, 0, 1, 15, -3, 0, -19, 0, 0, 0),
                (0, 0, 0, 0, 0, 0, 0, 0, 13, -9, 7, 1, -2, 0, 0),
                (0, 0, 0, 0, 0, -13, 0, -2, 13, 1, -3, -13, -13, 0, 0),
                (0, 0, 0, 0, 0, 0, 0, 6, -15, 3, -2, 8, -13, -13, 1),
                (0, 0, 0, 0, 0, 0, 0, -23, 0, 3, -7, -12, 6, 3, -7),
                (0, 0, 0, 0, 0, 0, 0, -20, 0, 0, -21, 12, -3, 0, 0),
                (0, 0, 0, 0, -31, 0, 0, 0, 18, -8, 0, 8, -1, -31, -31),
                (0, 0, 0, 0, 0, 0, 0, -8, -1, 4, 0, -9, 0, 7, -3)
                );
    constant parent : intArray2D(nTrees-1 downto 0)(nNodes-1 downto 0) := ((-1, 0, 0, 1, 1, 2, 2, 3, 3, 4, 4, 5, 5, 6, 6),
                (-1, 0, 0, 1, 1, 2, 2, 3, 3, 4, 4, 5, 5, 6, 6),
                (-1, 0, 0, 1, 1, 2, 2, 3, 3, 4, 4, 5, 5, 6, 6),
                (-1, 0, 0, 1, 1, 2, 2, 3, 3, 4, 4, 5, 5, 6, 6),
                (-1, 0, 0, 1, 1, 2, 2, 3, 3, 4, 4, 5, 5, 6, 6),
                (-1, 0, 0, 1, 1, 2, 2, 3, 3, 4, 4, 5, 5, 6, 6),
                (-1, 0, 0, 1, 1, 2, 2, 3, 3, 4, 4, 5, 5, 6, 6),
                (-1, 0, 0, 1, 1, 2, 2, 3, 3, 4, 4, 5, 5, 6, 6),
                (-1, 0, 0, 1, 1, 2, 2, 3, 3, 4, 4, 5, 5, 6, 6),
                (-1, 0, 0, 1, 1, 2, 2, 3, 3, 4, 4, 5, 5, 6, 6),
                (-1, 0, 0, 1, 1, 2, 2, 3, 3, 4, 4, 5, 5, 6, 6),
                (-1, 0, 0, 1, 1, 2, 2, 3, 3, 4, 4, 5, 5, 6, 6),
                (-1, 0, 0, 1, 1, 2, 2, 3, 3, 4, 4, 5, 5, 6, 6),
                (-1, 0, 0, 1, 1, 2, 2, 3, 3, 4, 4, 5, 5, 6, 6),
                (-1, 0, 0, 1, 1, 2, 2, 3, 3, 4, 4, 5, 5, 6, 6),
                (-1, 0, 0, 1, 1, 2, 2, 3, 3, 4, 4, 5, 5, 6, 6),
                (-1, 0, 0, 1, 1, 2, 2, 3, 3, 4, 4, 5, 5, 6, 6),
                (-1, 0, 0, 1, 1, 2, 2, 3, 3, 4, 4, 5, 5, 6, 6),
                (-1, 0, 0, 1, 1, 2, 2, 3, 3, 4, 4, 5, 5, 6, 6),
                (-1, 0, 0, 1, 1, 2, 2, 3, 3, 4, 4, 6, 6, 5, 5),
                (-1, 0, 0, 1, 1, 2, 2, 3, 3, 4, 4, 5, 5, 6, 6),
                (-1, 0, 0, 1, 1, 2, 2, 3, 3, 4, 4, 5, 5, 6, 6),
                (-1, 0, 0, 1, 1, 2, 2, 3, 3, 4, 4, 5, 5, 6, 6),
                (-1, 0, 0, 1, 1, 2, 2, 3, 3, 4, 4, 5, 5, 6, 6),
                (-1, 0, 0, 1, 1, 2, 2, 3, 3, 5, 5, 6, 6, 4, 4),
                (-1, 0, 0, 1, 1, 2, 2, 3, 3, 4, 4, 5, 5, 6, 6),
                (-1, 0, 0, 1, 1, 2, 2, 3, 3, 4, 4, 5, 5, 6, 6),
                (-1, 0, 0, 1, 1, 2, 2, 3, 3, 4, 4, 6, 6, 5, 5),
                (-1, 0, 0, 1, 1, 2, 2, 3, 3, 4, 4, 6, 6, 5, 5),
                (-1, 0, 0, 2, 2, 3, 3, 4, 4, 1, 1, 9, 9, 10, 10),
                (-1, 0, 0, 1, 1, 2, 2, 3, 3, 5, 5, 6, 6, 4, 4),
                (-1, 0, 0, 1, 1, 2, 2, 3, 3, 4, 4, 5, 5, 6, 6),
                (-1, 0, 0, 1, 1, 2, 2, 3, 3, 4, 4, 5, 5, 6, 6),
                (-1, 0, 0, 1, 1, 2, 2, 3, 3, 4, 4, 5, 5, 6, 6),
                (-1, 0, 0, 1, 1, 2, 2, 3, 3, 4, 4, 5, 5, 6, 6),
                (-1, 0, 0, 1, 1, 2, 2, 3, 3, 4, 4, 5, 5, 6, 6),
                (-1, 0, 0, 1, 1, 2, 2, 4, 4, 5, 5, 6, 6, 3, 3),
                (-1, 0, 0, 1, 1, 2, 2, 3, 3, 4, 4, 5, 5, 6, 6),
                (-1, 0, 0, 1, 1, 2, 2, 3, 3, 5, 5, 6, 6, 4, 4),
                (-1, 0, 0, 1, 1, 2, 2, 3, 3, 4, 4, 5, 5, 6, 6),
                (-1, 0, 0, 1, 1, 2, 2, 3, 3, 4, 4, 5, 5, 6, 6),
                (-1, 0, 0, 1, 1, 2, 2, 3, 3, 4, 4, 5, 5, 6, 6),
                (-1, 0, 0, 1, 1, 2, 2, 3, 3, 4, 4, 5, 5, 6, 6),
                (-1, 0, 0, 1, 1, 2, 2, 4, 4, 5, 5, 6, 6, 3, 3),
                (-1, 0, 0, 1, 1, 2, 2, 3, 3, 4, 4, 5, 5, 6, 6),
                (-1, 0, 0, 1, 1, 2, 2, 3, 3, 4, 4, 5, 5, 6, 6),
                (-1, 0, 0, 1, 1, 2, 2, 3, 3, 4, 4, 5, 5, 6, 6),
                (-1, 0, 0, 1, 1, 2, 2, 3, 3, 5, 5, 6, 6, 4, 4),
                (-1, 0, 0, 1, 1, 2, 2, 3, 3, 5, 5, 6, 6, 4, 4),
                (-1, 0, 0, 1, 1, 2, 2, 3, 3, 4, 4, 5, 5, 6, 6)
                );
    constant depth : intArray2D(nTrees-1 downto 0)(nNodes-1 downto 0) := ((0, 1, 1, 2, 2, 2, 2, 3, 3, 3, 3, 3, 3, 3, 3),
                (0, 1, 1, 2, 2, 2, 2, 3, 3, 3, 3, 3, 3, 3, 3),
                (0, 1, 1, 2, 2, 2, 2, 3, 3, 3, 3, 3, 3, 3, 3),
                (0, 1, 1, 2, 2, 2, 2, 3, 3, 3, 3, 3, 3, 3, 3),
                (0, 1, 1, 2, 2, 2, 2, 3, 3, 3, 3, 3, 3, 3, 3),
                (0, 1, 1, 2, 2, 2, 2, 3, 3, 3, 3, 3, 3, 3, 3),
                (0, 1, 1, 2, 2, 2, 2, 3, 3, 3, 3, 3, 3, 3, 3),
                (0, 1, 1, 2, 2, 2, 2, 3, 3, 3, 3, 3, 3, 3, 3),
                (0, 1, 1, 2, 2, 2, 2, 3, 3, 3, 3, 3, 3, 3, 3),
                (0, 1, 1, 2, 2, 2, 2, 3, 3, 3, 3, 3, 3, 3, 3),
                (0, 1, 1, 2, 2, 2, 2, 3, 3, 3, 3, 3, 3, 3, 3),
                (0, 1, 1, 2, 2, 2, 2, 3, 3, 3, 3, 3, 3, 3, 3),
                (0, 1, 1, 2, 2, 2, 2, 3, 3, 3, 3, 3, 3, 3, 3),
                (0, 1, 1, 2, 2, 2, 2, 3, 3, 3, 3, 3, 3, 3, 3),
                (0, 1, 1, 2, 2, 2, 2, 3, 3, 3, 3, 3, 3, 3, 3),
                (0, 1, 1, 2, 2, 2, 2, 3, 3, 3, 3, 3, 3, 3, 3),
                (0, 1, 1, 2, 2, 2, 2, 3, 3, 3, 3, 3, 3, 3, 3),
                (0, 1, 1, 2, 2, 2, 2, 3, 3, 3, 3, 3, 3, 3, 3),
                (0, 1, 1, 2, 2, 2, 2, 3, 3, 3, 3, 3, 3, 3, 3),
                (0, 1, 1, 2, 2, 2, 2, 3, 3, 3, 3, 3, 3, 3, 3),
                (0, 1, 1, 2, 2, 2, 2, 3, 3, 3, 3, 3, 3, 3, 3),
                (0, 1, 1, 2, 2, 2, 2, 3, 3, 3, 3, 3, 3, 3, 3),
                (0, 1, 1, 2, 2, 2, 2, 3, 3, 3, 3, 3, 3, 3, 3),
                (0, 1, 1, 2, 2, 2, 2, 3, 3, 3, 3, 3, 3, 3, 3),
                (0, 1, 1, 2, 2, 2, 2, 3, 3, 3, 3, 3, 3, 3, 3),
                (0, 1, 1, 2, 2, 2, 2, 3, 3, 3, 3, 3, 3, 3, 3),
                (0, 1, 1, 2, 2, 2, 2, 3, 3, 3, 3, 3, 3, 3, 3),
                (0, 1, 1, 2, 2, 2, 2, 3, 3, 3, 3, 3, 3, 3, 3),
                (0, 1, 1, 2, 2, 2, 2, 3, 3, 3, 3, 3, 3, 3, 3),
                (0, 1, 1, 2, 2, 3, 3, 3, 3, 2, 2, 3, 3, 3, 3),
                (0, 1, 1, 2, 2, 2, 2, 3, 3, 3, 3, 3, 3, 3, 3),
                (0, 1, 1, 2, 2, 2, 2, 3, 3, 3, 3, 3, 3, 3, 3),
                (0, 1, 1, 2, 2, 2, 2, 3, 3, 3, 3, 3, 3, 3, 3),
                (0, 1, 1, 2, 2, 2, 2, 3, 3, 3, 3, 3, 3, 3, 3),
                (0, 1, 1, 2, 2, 2, 2, 3, 3, 3, 3, 3, 3, 3, 3),
                (0, 1, 1, 2, 2, 2, 2, 3, 3, 3, 3, 3, 3, 3, 3),
                (0, 1, 1, 2, 2, 2, 2, 3, 3, 3, 3, 3, 3, 3, 3),
                (0, 1, 1, 2, 2, 2, 2, 3, 3, 3, 3, 3, 3, 3, 3),
                (0, 1, 1, 2, 2, 2, 2, 3, 3, 3, 3, 3, 3, 3, 3),
                (0, 1, 1, 2, 2, 2, 2, 3, 3, 3, 3, 3, 3, 3, 3),
                (0, 1, 1, 2, 2, 2, 2, 3, 3, 3, 3, 3, 3, 3, 3),
                (0, 1, 1, 2, 2, 2, 2, 3, 3, 3, 3, 3, 3, 3, 3),
                (0, 1, 1, 2, 2, 2, 2, 3, 3, 3, 3, 3, 3, 3, 3),
                (0, 1, 1, 2, 2, 2, 2, 3, 3, 3, 3, 3, 3, 3, 3),
                (0, 1, 1, 2, 2, 2, 2, 3, 3, 3, 3, 3, 3, 3, 3),
                (0, 1, 1, 2, 2, 2, 2, 3, 3, 3, 3, 3, 3, 3, 3),
                (0, 1, 1, 2, 2, 2, 2, 3, 3, 3, 3, 3, 3, 3, 3),
                (0, 1, 1, 2, 2, 2, 2, 3, 3, 3, 3, 3, 3, 3, 3),
                (0, 1, 1, 2, 2, 2, 2, 3, 3, 3, 3, 3, 3, 3, 3),
                (0, 1, 1, 2, 2, 2, 2, 3, 3, 3, 3, 3, 3, 3, 3)
                );
    constant iLeaf : intArray2D(nTrees-1 downto 0)(nLeaves-1 downto 0) := ((7, 8, 9, 10, 11, 12, 13, 14),
                (7, 8, 9, 10, 11, 12, 13, 14),
                (7, 8, 9, 10, 11, 12, 13, 14),
                (7, 8, 9, 10, 11, 12, 13, 14),
                (7, 8, 9, 10, 11, 12, 13, 14),
                (7, 8, 9, 10, 11, 12, 13, 14),
                (7, 8, 9, 10, 11, 12, 13, 14),
                (7, 8, 9, 10, 11, 12, 13, 14),
                (7, 8, 9, 10, 11, 12, 13, 14),
                (7, 8, 9, 10, 11, 12, 13, 14),
                (7, 8, 9, 10, 11, 12, 13, 14),
                (7, 8, 9, 10, 11, 12, 13, 14),
                (7, 8, 9, 10, 11, 12, 13, 14),
                (7, 8, 9, 10, 11, 12, 13, 14),
                (7, 8, 9, 10, 11, 12, 13, 14),
                (7, 8, 9, 10, 11, 12, 13, 14),
                (7, 8, 9, 10, 11, 12, 13, 14),
                (7, 8, 9, 10, 11, 12, 13, 14),
                (7, 8, 9, 10, 11, 12, 13, 14),
                (7, 8, 9, 10, 11, 12, 13, 14),
                (7, 8, 9, 10, 11, 12, 13, 14),
                (7, 8, 9, 10, 11, 12, 13, 14),
                (7, 8, 9, 10, 11, 12, 13, 14),
                (7, 8, 9, 10, 11, 12, 13, 14),
                (7, 8, 9, 10, 11, 12, 13, 14),
                (7, 8, 9, 10, 11, 12, 13, 14),
                (7, 8, 9, 10, 11, 12, 13, 14),
                (7, 8, 9, 10, 11, 12, 13, 14),
                (7, 8, 9, 10, 11, 12, 13, 14),
                (5, 6, 7, 8, 11, 12, 13, 14),
                (7, 8, 9, 10, 11, 12, 13, 14),
                (7, 8, 9, 10, 11, 12, 13, 14),
                (7, 8, 9, 10, 11, 12, 13, 14),
                (7, 8, 9, 10, 11, 12, 13, 14),
                (7, 8, 9, 10, 11, 12, 13, 14),
                (7, 8, 9, 10, 11, 12, 13, 14),
                (7, 8, 9, 10, 11, 12, 13, 14),
                (7, 8, 9, 10, 11, 12, 13, 14),
                (7, 8, 9, 10, 11, 12, 13, 14),
                (7, 8, 9, 10, 11, 12, 13, 14),
                (7, 8, 9, 10, 11, 12, 13, 14),
                (7, 8, 9, 10, 11, 12, 13, 14),
                (7, 8, 9, 10, 11, 12, 13, 14),
                (7, 8, 9, 10, 11, 12, 13, 14),
                (7, 8, 9, 10, 11, 12, 13, 14),
                (7, 8, 9, 10, 11, 12, 13, 14),
                (7, 8, 9, 10, 11, 12, 13, 14),
                (7, 8, 9, 10, 11, 12, 13, 14),
                (7, 8, 9, 10, 11, 12, 13, 14),
                (7, 8, 9, 10, 11, 12, 13, 14)
                );
    constant value : tyArray2D(nTrees-1 downto 0)(nNodes-1 downto 0) := to_tyArray2D(value_int);
      constant threshold : txArray2D(nTrees-1 downto 0)(nNodes-1 downto 0) := to_txArray2D(threshold_int);
end Arrays0;