library ieee;
use ieee.std_logic_1164.all;
use ieee.std_logic_misc.all;
use ieee.numeric_std.all;

package TanLROM is
    type intArray is array(natural range <>) of integer;
    type intArray2D is array(natural range <>) of intArray;

    constant Phi_shift : intArray(0 TO 17) := (
        (0),(0),
        (86),(86),
        (172),(172),
        (258),(258),
        (344),(344),
        (430),(430),
        (516),(516),
        (602),(602),
        (688),(688));
 
     
    constant TanLLUT : intArray2D(0 to 127)(0 to 6) := (
        (2,342,559,704,810,894,964),
(5,344,560,704,811,895,964),
(7,346,561,705,812,896,965),
(10,348,562,707,813,896,965),
(13,350,565,708,813,897,966),
(15,353,566,709,814,897,966),
(21,355,567,709,815,898,967),
(23,357,568,710,815,898,968),
(26,359,569,711,816,899,968),
(29,360,571,712,817,900,968),
(31,362,572,713,818,901,969),
(34,364,574,714,818,901,969),
(37,368,575,715,819,902,970),
(42,369,576,716,820,902,970),
(44,371,577,717,820,903,971),
(47,373,579,718,821,904,971),
(50,375,580,718,822,904,972),
(52,376,581,720,823,905,972),
(55,380,583,721,823,905,973),
(60,382,584,722,824,906,973),
(63,383,585,722,825,906,974),
(65,385,586,723,825,907,974),
(68,387,587,724,827,908,975),
(71,389,589,726,827,908,975),
(73,390,591,726,828,909,976),
(76,394,592,727,828,909,976),
(81,395,593,728,829,910,976),
(84,397,594,729,830,910,977),
(86,399,595,729,830,911,978),
(89,400,596,730,831,912,978),
(91,402,597,732,832,912,979),
(94,404,599,733,833,913,979),
(96,407,601,733,833,913,979),
(102,409,602,734,834,914,980),
(104,410,603,735,834,914,981),
(107,412,604,736,835,915,981),
(109,414,605,737,836,916,981),
(112,415,607,738,837,916,982),
(114,418,608,739,837,917,982),
(119,420,609,740,838,917,983),
(122,422,610,740,839,918,984),
(124,423,611,741,839,918,984),
(127,425,612,742,840,919,984),
(129,426,613,743,841,919,985),
(132,428,615,744,842,920,985),
(134,431,616,745,842,920,986),
(139,433,617,746,843,921,986),
(142,434,618,746,843,921,987),
(144,436,619,747,844,922,987),
(147,437,620,748,845,923,988),
(149,439,621,749,846,923,988),
(152,440,623,750,846,924,988),
(154,443,624,751,847,924,989),
(159,445,625,752,848,925,989),
(162,447,626,752,848,926,990),
(164,448,628,753,849,926,991),
(166,450,629,755,850,927,991),
(169,451,631,755,850,927,991),
(171,454,632,756,851,928,992),
(176,456,633,757,852,928,992),
(178,457,633,757,852,929,993),
(181,458,634,758,853,930,993),
(183,460,635,759,854,930,994),
(186,461,636,760,854,930,994),
(188,463,638,761,855,931,995),
(190,466,639,762,856,931,995),
(195,467,640,763,856,932,995),
(197,469,641,763,857,932,996),
(200,470,642,764,857,933,997),
(202,472,643,765,858,934,997),
(204,473,644,766,859,934,997),
(207,474,646,767,860,935,998),
(211,477,647,768,860,935,998),
(213,479,648,768,861,936,999),
(216,480,649,769,861,937,999),
(218,482,650,770,862,937,1000),
(220,483,651,771,863,938,1000),
(223,484,653,772,864,938,1001),
(225,487,654,773,864,938,1001),
(229,489,655,773,865,939,1001),
(232,490,656,774,865,939,1002),
(234,491,657,775,866,940,1003),
(236,493,658,775,867,941,1003),
(238,494,658,777,867,941,1003),
(240,495,660,777,868,942,1004),
(243,498,661,778,869,942,1004),
(247,499,662,779,869,943,1004),
(249,501,663,780,870,943,1005),
(251,502,664,780,870,944,1006),
(254,504,665,781,871,944,1006),
(256,505,667,782,872,945,1006),
(258,508,668,783,872,945,1007),
(262,509,669,784,873,946,1007),
(264,510,670,784,874,946,1008),
(266,511,670,785,874,947,1008),
(269,513,671,786,875,948,1009),
(271,514,672,787,876,948,1009),
(273,515,674,788,876,949,1010),
(275,518,675,788,877,949,1010),
(279,519,676,789,877,949,1010),
(281,521,677,790,878,950,1011),
(283,522,678,790,878,951,1011),
(285,523,679,791,880,951,1012),
(287,524,679,792,880,952,1012),
(289,526,681,793,881,952,1013),
(291,528,682,794,881,953,1013),
(295,530,683,795,882,953,1013),
(297,531,684,795,882,953,1014),
(299,532,685,796,883,954,1015),
(301,533,686,797,884,955,1015),
(303,535,687,798,884,955,1015),
(305,537,688,798,885,956,1016),
(309,538,689,799,885,956,1016),
(311,540,690,800,886,957,1017),
(313,541,691,800,886,957,1017),
(315,542,692,801,888,958,1018),
(317,543,693,802,888,958,1018),
(319,544,694,803,889,959,1018),
(321,547,695,804,889,959,1019),
(325,548,696,804,890,960,1019),
(327,549,697,805,890,960,1020),
(329,551,698,806,891,961,1020),
(331,552,698,806,892,961,1021),
(333,553,699,808,892,962,1021),
(335,554,701,808,893,962,1021),
(336,557,702,809,893,963,1022),
(340,558,703,810,894,963,1022),
(0,0,0,0,0,0,0)        
);


end TanLROM; 