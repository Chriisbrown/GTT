../../../../RuflCore/firmware/hdl/ReuseableElements/PkgArrayTypes.vhd