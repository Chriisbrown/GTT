library ieee;
use ieee.std_logic_1164.all;
use ieee.std_logic_misc.all;
use ieee.numeric_std.all;

package TanLROM is
    type intArray is array(natural range <>) of integer;
    type intArray2D is array(natural range <>) of intArray;

    constant Phi_shift : intArray(0 TO 17) := (
        (0),(0),
      (696),(696),
     (1392),(1392),
     (2088),(2088),
     (2784),(2784),
     (3480),(3480),
     (4176),(4176),
     (4872),(4872),
     (5568),(5568));
     
    constant TanLLUT : intArray2D(0 to 4095)(0 to 7) := (
        (32769,43691,50658,55303,58727,61425,63647,65535),
        (32771,43693,50659,55304,58728,61425,63648,0),
        (32774,43695,50661,55305,58728,61426,63648,0),
        (32778,43697,50662,55306,58729,61426,63649,0),
        (32781,43699,50664,55307,58729,61427,63649,0),
        (32783,43701,50665,55308,58730,61428,63650,0),
        (32786,43704,50667,55309,58731,61428,63650,0),
        (32790,43706,50668,55310,58732,61429,63651,0),
        (32793,43708,50669,55311,58733,61430,63651,0),
        (32795,43710,50671,55312,58733,61430,63652,0),
        (32799,43712,50672,55313,58734,61431,63652,0),
        (32802,43714,50673,55313,58735,61431,63653,0),
        (32805,43716,50674,55315,58736,61432,63653,0),
        (32807,43719,50676,55316,58736,61432,63654,0),
        (32811,43721,50677,55316,58737,61433,63654,0),
        (32814,43723,50678,55317,58738,61434,63655,0),
        (32816,43724,50680,55318,58738,61434,63655,0),
        (32820,43727,50681,55319,58739,61435,63656,0),
        (32823,43729,50683,55320,58740,61436,63656,0),
        (32826,43731,50684,55321,58741,61436,63657,0),
        (32828,43734,50686,55322,58741,61437,63657,0),
        (32832,43736,50687,55323,58742,61437,63658,0),
        (32835,43738,50688,55324,58743,61438,63658,0),
        (32838,43739,50690,55325,58744,61438,63659,0),
        (32842,43742,50691,55326,58744,61439,63659,0),
        (32844,43744,50692,55327,58745,61440,63660,0),
        (32847,43746,50693,55328,58746,61440,63660,0),
        (32850,43749,50695,55329,58746,61441,63661,0),
        (32854,43751,50696,55330,58747,61441,63661,0),
        (32856,43752,50697,55331,58748,61442,63662,0),
        (32859,43754,50699,55332,58749,61443,63662,0),
        (32863,43757,50700,55333,58749,61443,63663,0),
        (32865,43759,50701,55334,58750,61444,63663,0),
        (32868,43761,50703,55335,58751,61444,63664,0),
        (32871,43764,50704,55336,58752,61445,63664,0),
        (32875,43766,50706,55336,58752,61445,63665,0),
        (32877,43767,50707,55337,58753,61446,63665,0),
        (32880,43769,50709,55339,58754,61447,63666,0),
        (32884,43772,50710,55339,58754,61447,63666,0),
        (32887,43774,50711,55340,58755,61448,63667,0),
        (32889,43776,50712,55341,58756,61449,63667,0),
        (32892,43779,50714,55342,58757,61449,63668,0),
        (32896,43780,50715,55343,58757,61450,63668,0),
        (32899,43782,50716,55344,58758,61450,63669,0),
        (32901,43784,50718,55345,58759,61451,63669,0),
        (32905,43787,50719,55346,58760,61451,63670,0),
        (32908,43789,50720,55347,58760,61452,63670,0),
        (32910,43791,50721,55348,58761,61453,63671,0),
        (32913,43793,50723,55349,58762,61453,63671,0),
        (32917,43795,50724,55350,58762,61454,63672,0),
        (32920,43797,50726,55351,58763,61454,63672,0),
        (32922,43799,50727,55352,58764,61455,63673,0),
        (32926,43802,50729,55353,58765,61456,63673,0),
        (32929,43804,50730,55354,58765,61456,63674,0),
        (32932,43806,50731,55355,58766,61457,63674,0),
        (32934,43808,50733,55356,58767,61457,63675,0),
        (32938,43810,50734,55356,58768,61458,63675,0),
        (32941,43812,50735,55357,58769,61459,63676,0),
        (32944,43814,50737,55359,58769,61459,63676,0),
        (32948,43817,50738,55359,58770,61460,63676,0),
        (32950,43819,50739,55360,58770,61460,63677,0),
        (32953,43820,50740,55361,58771,61461,63678,0),
        (32955,43823,50742,55362,58772,61461,63678,0),
        (32959,43825,50743,55363,58773,61462,63679,0),
        (32962,43827,50744,55364,58774,61463,63679,0),
        (32965,43829,50746,55365,58774,61463,63680,0),
        (32969,43832,50747,55366,58775,61464,63680,0),
        (32971,43833,50749,55367,58776,61465,63681,0),
        (32974,43835,50750,55368,58777,61465,63681,0),
        (32977,43838,50752,55369,58777,61466,63681,0),
        (32981,43840,50753,55370,58778,61466,63682,0),
        (32983,43842,50754,55371,58779,61467,63683,0),
        (32986,43844,50756,55372,58779,61467,63683,0),
        (32990,43846,50757,55373,58780,61468,63683,0),
        (32993,43848,50758,55374,58781,61469,63684,0),
        (32995,43850,50759,55375,58782,61469,63685,0),
        (32998,43853,50761,55376,58782,61470,63685,0),
        (33002,43855,50762,55376,58783,61470,63686,0),
        (33004,43857,50763,55377,58784,61471,63686,0),
        (33007,43858,50765,55379,58785,61472,63686,0),
        (33011,43861,50766,55379,58785,61472,63687,0),
        (33014,43863,50767,55380,58786,61473,63688,0),
        (33016,43865,50769,55381,58787,61473,63688,0),
        (33019,43868,50770,55382,58787,61474,63688,0),
        (33023,43870,50771,55383,58788,61474,63689,0),
        (33026,43871,50773,55384,58789,61475,63689,0),
        (33028,43873,50774,55385,58790,61476,63690,0),
        (33032,43876,50776,55386,58790,61476,63690,0),
        (33035,43878,50777,55387,58791,61477,63691,0),
        (33038,43880,50778,55388,58792,61478,63691,0),
        (33040,43883,50780,55389,58793,61478,63692,0),
        (33044,43884,50781,55390,58793,61479,63693,0),
        (33047,43886,50782,55391,58794,61479,63693,0),
        (33049,43888,50784,55392,58795,61480,63693,0),
        (33053,43891,50785,55393,58795,61480,63694,0),
        (33056,43893,50786,55394,58796,61481,63694,0),
        (33059,43895,50787,55395,58797,61482,63695,0),
        (33061,43897,50789,55396,58798,61482,63695,0),
        (33065,43899,50790,55396,58798,61483,63696,0),
        (33068,43901,50791,55397,58799,61483,63696,0),
        (33071,43903,50793,55399,58800,61484,63697,0),
        (33075,43906,50794,55399,58800,61484,63697,0),
        (33077,43908,50796,55400,58801,61485,63698,0),
        (33080,43909,50797,55401,58802,61486,63698,0),
        (33083,43912,50798,55402,58803,61486,63699,0),
        (33086,43914,50800,55403,58803,61487,63699,0),
        (33089,43916,50801,55404,58804,61488,63700,0),
        (33092,43918,50803,55405,58805,61488,63700,0),
        (33096,43920,50804,55406,58806,61489,63701,0),
        (33098,43922,50805,55407,58806,61489,63701,0),
        (33101,43924,50806,55408,58807,61490,63702,0),
        (33104,43927,50808,55409,58808,61490,63702,0),
        (33108,43929,50809,55410,58808,61491,63703,0),
        (33110,43931,50810,55411,58809,61492,63703,0),
        (33113,43932,50812,55412,58810,61492,63704,0),
        (33117,43935,50813,55413,58811,61493,63704,0),
        (33120,43937,50814,55413,58811,61494,63705,0),
        (33122,43939,50815,55415,58812,61494,63705,0),
        (33125,43942,50817,55416,58813,61495,63706,0),
        (33129,43944,50818,55416,58814,61495,63706,0),
        (33131,43945,50820,55417,58815,61496,63707,0),
        (33134,43947,50821,55418,58815,61496,63707,0),
        (33138,43950,50822,55419,58816,61497,63708,0),
        (33141,43952,50824,55420,58816,61498,63708,0),
        (33143,43954,50825,55421,58817,61498,63709,0),
        (33146,43956,50827,55422,58818,61499,63709,0),
        (33150,43958,50828,55423,58819,61499,63710,0),
        (33153,43960,50829,55424,58820,61500,63710,0),
        (33155,43962,50831,55425,58820,61501,63711,0),
        (33159,43965,50832,55426,58821,61501,63711,0),
        (33162,43967,50833,55427,58822,61502,63712,0),
        (33165,43968,50834,55428,58822,61502,63712,0),
        (33167,43971,50836,55429,58823,61503,63713,0),
        (33171,43973,50837,55430,58824,61503,63713,0),
        (33174,43975,50838,55430,58825,61504,63714,0),
        (33176,43977,50840,55432,58825,61505,63714,0),
        (33180,43979,50841,55433,58826,61505,63715,0),
        (33183,43981,50842,55433,58827,61506,63715,0),
        (33186,43983,50844,55435,58828,61506,63716,0),
        (33188,43986,50845,55435,58828,61507,63716,0),
        (33192,43988,50846,55436,58829,61507,63717,0),
        (33195,43990,50848,55437,58830,61508,63717,0),
        (33198,43991,50849,55438,58830,61509,63718,0),
        (33202,43994,50851,55439,58831,61509,63718,0),
        (33204,43996,50852,55440,58832,61510,63719,0),
        (33207,43998,50853,55441,58833,61511,63719,0),
        (33210,44001,50855,55442,58833,61511,63720,0),
        (33213,44002,50856,55443,58834,61512,63720,0),
        (33216,44004,50857,55444,58835,61512,63721,0),
        (33219,44006,50859,55445,58836,61513,63721,0),
        (33223,44009,50860,55446,58836,61513,63722,0),
        (33225,44011,50861,55447,58837,61514,63722,0),
        (33228,44013,50862,55448,58838,61515,63723,0),
        (33231,44015,50864,55449,58838,61515,63723,0),
        (33235,44017,50865,55450,58839,61516,63724,0),
        (33237,44019,50866,55450,58840,61516,63724,0),
        (33240,44021,50868,55452,58841,61517,63725,0),
        (33244,44024,50869,55452,58841,61518,63725,0),
        (33247,44025,50870,55453,58842,61518,63726,0),
        (33249,44027,50872,55454,58843,61519,63726,0),
        (33252,44030,50873,55455,58844,61519,63727,0),
        (33256,44032,50874,55456,58844,61520,63727,0),
        (33258,44034,50876,55457,58845,61521,63728,0),
        (33261,44036,50877,55458,58846,61521,63728,0),
        (33265,44038,50879,55459,58846,61522,63728,0),
        (33268,44040,50880,55460,58847,61522,63729,0),
        (33270,44042,50881,55461,58848,61523,63730,0),
        (33273,44045,50883,55462,58849,61523,63730,0),
        (33277,44047,50884,55463,58849,61524,63731,0),
        (33280,44048,50885,55464,58850,61525,63731,0),
        (33282,44050,50887,55465,58851,61525,63732,0),
        (33286,44053,50888,55466,58851,61526,63732,0),
        (33289,44055,50889,55466,58852,61527,63733,0),
        (33292,44057,50890,55468,58853,61527,63733,0),
        (33294,44059,50892,55469,58854,61528,63733,0),
        (33298,44061,50893,55469,58854,61528,63734,0),
        (33301,44063,50894,55470,58855,61529,63735,0),
        (33303,44065,50896,55471,58856,61529,63735,0),
        (33307,44068,50897,55472,58857,61530,63735,0),
        (33310,44069,50898,55473,58857,61531,63736,0),
        (33313,44071,50899,55474,58858,61531,63736,0),
        (33315,44074,50901,55475,58859,61532,63737,0),
        (33319,44076,50902,55476,58859,61532,63738,0),
        (33322,44078,50904,55477,58860,61533,63738,0),
        (33325,44080,50905,55478,58861,61533,63738,0),
        (33329,44082,50906,55479,58862,61534,63739,0),
        (33331,44084,50908,55480,58862,61535,63739,0),
        (33334,44086,50909,55481,58863,61535,63740,0),
        (33336,44089,50911,55482,58864,61536,63740,0),
        (33340,44091,50912,55483,58864,61536,63741,0),
        (33343,44092,50913,55483,58865,61537,63741,0),
        (33346,44094,50915,55485,58866,61538,63742,0),
        (33350,44097,50916,55485,58867,61538,63742,0),
        (33352,44099,50917,55486,58867,61539,63743,0),
        (33355,44101,50918,55488,58868,61539,63743,0),
        (33358,44103,50920,55488,58869,61540,63744,0),
        (33362,44105,50921,55489,58870,61540,63744,0),
        (33364,44107,50922,55490,58871,61541,63745,0),
        (33367,44109,50924,55491,58871,61542,63745,0),
        (33371,44112,50925,55492,58872,61542,63746,0),
        (33374,44113,50926,55493,58872,61543,63746,0),
        (33376,44115,50927,55494,58873,61544,63747,0),
        (33379,44118,50929,55495,58874,61544,63747,0),
        (33383,44120,50930,55496,58875,61545,63748,0),
        (33385,44122,50931,55497,58876,61545,63748,0),
        (33388,44123,50933,55498,58876,61546,63749,0),
        (33392,44126,50934,55499,58877,61546,63749,0),
        (33395,44128,50936,55499,58878,61547,63750,0),
        (33397,44130,50937,55501,58878,61548,63750,0),
        (33400,44133,50938,55502,58879,61548,63751,0),
        (33404,44134,50940,55502,58880,61549,63751,0),
        (33407,44136,50941,55503,58881,61549,63752,0),
        (33409,44138,50942,55504,58881,61550,63752,0),
        (33413,44141,50944,55505,58882,61550,63753,0),
        (33416,44143,50945,55506,58883,61551,63753,0),
        (33418,44144,50946,55507,58884,61552,63754,0),
        (33421,44147,50948,55508,58884,61552,63754,0),
        (33425,44149,50949,55509,58885,61553,63755,0),
        (33428,44151,50950,55510,58886,61554,63755,0),
        (33430,44153,50952,55511,58886,61554,63756,0),
        (33434,44155,50953,55512,58887,61555,63756,0),
        (33437,44157,50954,55513,58888,61555,63757,0),
        (33440,44159,50955,55514,58889,61556,63757,0),
        (33442,44162,50957,55515,58889,61556,63758,0),
        (33446,44164,50958,55516,58890,61557,63758,0),
        (33449,44165,50959,55516,58891,61558,63759,0),
        (33452,44167,50961,55518,58891,61558,63759,0),
        (33455,44170,50962,55518,58892,61559,63760,0),
        (33458,44172,50963,55519,58893,61559,63760,0),
        (33461,44174,50964,55521,58894,61560,63761,0),
        (33463,44176,50966,55521,58894,61560,63761,0),
        (33467,44178,50967,55522,58895,61561,63762,0),
        (33470,44180,50969,55523,58896,61562,63762,0),
        (33473,44182,50970,55524,58897,61562,63763,0),
        (33477,44184,50971,55525,58897,61563,63763,0),
        (33479,44186,50973,55526,58898,61564,63764,0),
        (33482,44188,50974,55527,58899,61564,63764,0),
        (33485,44191,50975,55528,58899,61565,63765,0),
        (33489,44193,50977,55529,58900,61565,63765,0),
        (33491,44194,50978,55530,58901,61566,63766,0),
        (33494,44196,50980,55531,58902,61566,63766,0),
        (33498,44199,50981,55532,58902,61567,63766,0),
        (33500,44201,50982,55532,58903,61568,63767,0),
        (33503,44203,50983,55534,58904,61568,63768,0),
        (33506,44205,50985,55535,58904,61569,63768,0),
        (33510,44207,50986,55535,58905,61569,63769,0),
        (33512,44209,50987,55536,58906,61570,63769,0),
        (33515,44211,50989,55537,58907,61570,63769,0),
        (33519,44214,50990,55538,58907,61571,63770,0),
        (33522,44215,50991,55539,58908,61572,63771,0),
        (33524,44217,50992,55540,58909,61572,63771,0),
        (33527,44220,50994,55541,58910,61573,63771,0),
        (33531,44222,50995,55542,58910,61573,63772,0),
        (33533,44224,50996,55543,58911,61574,63773,0),
        (33536,44225,50998,55544,58912,61575,63773,0),
        (33540,44228,50999,55545,58912,61575,63773,0),
        (33543,44230,51000,55546,58913,61576,63774,0),
        (33545,44232,51001,55547,58914,61576,63774,0),
        (33548,44234,51003,55548,58915,61577,63775,0),
        (33552,44236,51004,55548,58915,61577,63776,0),
        (33555,44238,51006,55549,58916,61578,63776,0),
        (33557,44240,51007,55551,58917,61579,63776,0),
        (33561,44243,51008,55551,58917,61579,63777,0),
        (33564,44244,51010,55552,58918,61580,63777,0),
        (33566,44246,51011,55553,58919,61581,63778,0),
        (33569,44249,51012,55554,58920,61581,63778,0),
        (33573,44251,51014,55555,58920,61582,63779,0),
        (33576,44253,51015,55556,58921,61582,63779,0),
        (33578,44254,51016,55557,58922,61583,63780,0),
        (33582,44257,51018,55558,58922,61583,63780,0),
        (33585,44259,51019,55559,58923,61584,63781,0),
        (33588,44261,51020,55560,58924,61585,63781,0),
        (33590,44263,51022,55561,58925,61585,63782,0),
        (33594,44265,51023,55562,58925,61586,63782,0),
        (33597,44267,51024,55563,58926,61586,63783,0),
        (33599,44270,51026,55564,58927,61587,63783,0),
        (33603,44272,51027,55564,58928,61587,63784,0),
        (33606,44273,51028,55565,58928,61588,63784,0),
        (33609,44275,51030,55567,58929,61589,63785,0),
        (33613,44278,51031,55567,58930,61589,63785,0),
        (33615,44280,51032,55568,58930,61590,63786,0),
        (33618,44282,51033,55569,58931,61590,63786,0),
        (33621,44284,51035,55570,58932,61591,63787,0),
        (33625,44286,51036,55571,58933,61592,63787,0),
        (33627,44288,51037,55572,58934,61592,63788,0),
        (33630,44290,51039,55573,58934,61593,63788,0),
        (33634,44292,51040,55574,58935,61593,63789,0),
        (33636,44294,51041,55575,58935,61594,63789,0),
        (33639,44296,51042,55576,58936,61595,63790,0),
        (33642,44299,51044,55577,58937,61595,63790,0),
        (33646,44300,51045,55578,58938,61596,63791,0),
        (33648,44302,51046,55578,58939,61596,63791,0),
        (33651,44304,51048,55580,58939,61597,63792,0),
        (33655,44307,51049,55580,58940,61597,63792,0),
        (33658,44309,51050,55581,58940,61598,63793,0),
        (33660,44310,51052,55583,58941,61599,63793,0),
        (33663,44313,51053,55583,58942,61599,63794,0),
        (33667,44315,51055,55584,58943,61600,63794,0),
        (33669,44317,51056,55585,58944,61600,63795,0),
        (33672,44319,51057,55586,58944,61601,63795,0),
        (33676,44321,51059,55587,58945,61602,63796,0),
        (33679,44323,51060,55588,58946,61602,63796,0),
        (33681,44325,51061,55589,58946,61603,63797,0),
        (33684,44328,51063,55590,58947,61603,63797,0),
        (33688,44329,51064,55591,58948,61604,63798,0),
        (33691,44331,51065,55592,58949,61605,63798,0),
        (33693,44333,51067,55593,58949,61605,63799,0),
        (33697,44336,51068,55594,58950,61606,63799,0),
        (33700,44337,51069,55594,58951,61606,63800,0),
        (33702,44339,51070,55596,58952,61607,63800,0),
        (33705,44342,51072,55596,58952,61607,63800,0),
        (33709,44344,51073,55597,58953,61608,63801,0),
        (33712,44346,51074,55598,58954,61609,63802,0),
        (33714,44347,51076,55599,58954,61609,63802,0),
        (33718,44350,51077,55600,58955,61610,63802,0),
        (33721,44352,51078,55601,58956,61610,63803,0),
        (33724,44354,51079,55602,58957,61611,63803,0),
        (33726,44356,51081,55603,58957,61611,63804,0),
        (33730,44358,51082,55604,58958,61612,63805,0),
        (33733,44360,51083,55605,58959,61613,63805,0),
        (33735,44362,51085,55606,58959,61613,63805,0),
        (33739,44365,51086,55607,58960,61614,63806,0),
        (33742,44366,51087,55607,58961,61615,63806,0),
        (33745,44368,51088,55609,58962,61615,63807,0),
        (33747,44371,51090,55610,58962,61616,63807,0),
        (33751,44373,51091,55610,58963,61616,63808,0),
        (33754,44374,51092,55611,58964,61617,63808,0),
        (33757,44376,51094,55612,58964,61617,63809,0),
        (33761,44379,51095,55613,58965,61618,63809,0),
        (33763,44381,51096,55614,58966,61619,63810,0),
        (33766,44382,51098,55615,58967,61619,63810,0),
        (33768,44385,51099,55616,58967,61620,63811,0),
        (33772,44387,51100,55617,58968,61620,63811,0),
        (33775,44389,51102,55618,58969,61621,63812,0),
        (33778,44391,51103,55619,58969,61621,63812,0),
        (33782,44393,51104,55620,58970,61622,63813,0),
        (33784,44395,51106,55621,58971,61623,63813,0),
        (33787,44397,51107,55622,58972,61623,63814,0),
        (33790,44400,51108,55623,58972,61624,63814,0),
        (33794,44401,51110,55623,58973,61624,63815,0),
        (33796,44403,51111,55624,58974,61625,63815,0),
        (33799,44405,51112,55625,58975,61626,63816,0),
        (33803,44408,51114,55626,58975,61626,63816,0),
        (33805,44409,51115,55627,58976,61627,63817,0),
        (33808,44411,51116,55628,58977,61627,63817,0),
        (33811,44414,51118,55629,58977,61628,63818,0),
        (33815,44416,51119,55630,58978,61628,63818,0),
        (33817,44418,51120,55631,58979,61629,63819,0),
        (33820,44419,51122,55632,58980,61630,63819,0),
        (33824,44422,51123,55633,58980,61630,63820,0),
        (33826,44424,51124,55634,58981,61631,63820,0),
        (33829,44426,51125,55635,58982,61631,63821,0),
        (33832,44428,51127,55636,58982,61632,63821,0),
        (33836,44430,51128,55636,58983,61632,63822,0),
        (33838,44432,51129,55637,58984,61633,63822,0),
        (33841,44434,51131,55639,58985,61634,63823,0),
        (33845,44436,51132,55639,58985,61634,63823,0),
        (33848,44438,51133,55640,58986,61635,63824,0),
        (33850,44440,51134,55641,58987,61636,63824,0),
        (33853,44443,51136,55642,58987,61636,63825,0),
        (33857,44444,51137,55643,58988,61637,63825,0),
        (33859,44446,51138,55644,58989,61637,63826,0),
        (33862,44448,51140,55645,58990,61638,63826,0),
        (33866,44451,51141,55646,58990,61638,63826,0),
        (33869,44452,51142,55647,58991,61639,63827,0),
        (33871,44454,51143,55648,58992,61640,63828,0),
        (33874,44457,51145,55649,58992,61640,63828,0),
        (33878,44459,51146,55650,58993,61641,63829,0),
        (33881,44461,51147,55650,58994,61641,63829,0),
        (33883,44462,51149,55652,58995,61642,63829,0),
        (33887,44465,51150,55652,58995,61642,63830,0),
        (33890,44467,51151,55653,58996,61643,63831,0),
        (33892,44469,51153,55654,58997,61644,63831,0),
        (33895,44471,51154,55655,58997,61644,63831,0),
        (33899,44473,51155,55656,58998,61645,63832,0),
        (33902,44475,51157,55657,58999,61645,63832,0),
        (33904,44477,51158,55658,59000,61646,63833,0),
        (33908,44479,51159,55659,59000,61646,63833,0),
        (33911,44481,51161,55660,59001,61647,63834,0),
        (33914,44483,51162,55661,59002,61648,63834,0),
        (33916,44486,51163,55662,59003,61648,63835,0),
        (33920,44487,51165,55663,59003,61649,63835,0),
        (33923,44489,51166,55663,59004,61650,63836,0),
        (33925,44491,51167,55665,59005,61650,63836,0),
        (33929,44494,51169,55665,59005,61651,63837,0),
        (33932,44495,51170,55666,59006,61651,63837,0),
        (33935,44497,51171,55667,59007,61652,63838,0),
        (33937,44500,51172,55668,59008,61652,63838,0),
        (33941,44502,51174,55669,59008,61653,63839,0),
        (33944,44503,51175,55670,59009,61654,63839,0),
        (33946,44505,51176,55671,59010,61654,63840,0),
        (33950,44508,51178,55672,59010,61655,63840,0),
        (33953,44510,51179,55673,59011,61655,63841,0),
        (33956,44511,51180,55674,59012,61656,63841,0),
        (33958,44514,51182,55675,59013,61656,63842,0),
        (33962,44516,51183,55676,59013,61657,63842,0),
        (33965,44518,51184,55676,59014,61658,63843,0),
        (33968,44519,51186,55678,59015,61658,63843,0),
        (33971,44522,51187,55678,59015,61659,63844,0),
        (33974,44524,51188,55679,59016,61659,63844,0),
        (33977,44526,51189,55680,59017,61660,63845,0),
        (33979,44528,51191,55681,59018,61661,63845,0),
        (33983,44530,51192,55682,59018,61661,63846,0),
        (33986,44532,51193,55683,59019,61662,63846,0),
        (33989,44534,51195,55684,59020,61662,63847,0),
        (33993,44536,51196,55685,59020,61663,63847,0),
        (33995,44538,51197,55686,59021,61664,63848,0),
        (33998,44540,51198,55687,59022,61664,63848,0),
        (34000,44543,51200,55688,59023,61665,63849,0),
        (34004,44544,51201,55689,59023,61665,63849,0),
        (34007,44546,51202,55689,59024,61666,63850,0),
        (34010,44548,51204,55691,59025,61666,63850,0),
        (34014,44551,51205,55691,59025,61667,63850,0),
        (34016,44552,51206,55692,59026,61668,63851,0),
        (34019,44554,51207,55693,59027,61668,63852,0),
        (34022,44557,51209,55694,59028,61669,63852,0),
        (34025,44559,51210,55695,59028,61669,63853,0),
        (34028,44560,51211,55696,59029,61670,63853,0),
        (34031,44562,51213,55697,59030,61670,63853,0),
        (34035,44565,51214,55698,59030,61671,63854,0),
        (34037,44567,51215,55699,59031,61672,63855,0),
        (34040,44568,51216,55700,59032,61672,63855,0),
        (34043,44571,51218,55701,59033,61673,63855,0),
        (34047,44573,51219,55702,59033,61673,63856,0),
        (34049,44575,51220,55702,59034,61674,63856,0),
        (34052,44576,51222,55704,59035,61675,63857,0),
        (34056,44579,51223,55704,59035,61675,63857,0),
        (34058,44581,51224,55705,59036,61676,63858,0),
        (34061,44583,51225,55706,59037,61676,63858,0),
        (34064,44585,51227,55707,59038,61677,63859,0),
        (34068,44587,51228,55708,59038,61677,63859,0),
        (34070,44589,51229,55709,59039,61678,63860,0),
        (34073,44591,51231,55710,59040,61679,63860,0),
        (34077,44593,51232,55711,59040,61679,63861,0),
        (34079,44595,51233,55712,59041,61680,63861,0),
        (34082,44597,51235,55713,59042,61680,63862,0),
        (34085,44600,51236,55714,59043,61681,63862,0),
        (34089,44601,51237,55715,59043,61681,63863,0),
        (34091,44603,51238,55715,59044,61682,63863,0),
        (34094,44605,51240,55717,59045,61683,63864,0),
        (34098,44608,51241,55717,59045,61683,63864,0),
        (34101,44609,51242,55718,59046,61684,63865,0),
        (34103,44611,51244,55719,59047,61684,63865,0),
        (34106,44614,51245,55720,59048,61685,63866,0),
        (34110,44616,51246,55721,59048,61685,63866,0),
        (34112,44617,51248,55722,59049,61686,63867,0),
        (34115,44619,51249,55723,59050,61687,63867,0),
        (34119,44622,51250,55724,59051,61687,63868,0),
        (34122,44624,51252,55725,59051,61688,63868,0),
        (34124,44625,51253,55726,59052,61689,63869,0),
        (34127,44628,51254,55727,59053,61689,63869,0),
        (34131,44630,51256,55728,59053,61690,63870,0),
        (34133,44631,51257,55728,59054,61690,63870,0),
        (34136,44633,51258,55730,59055,61691,63871,0),
        (34140,44636,51259,55730,59056,61691,63871,0),
        (34143,44638,51261,55731,59056,61692,63872,0),
        (34145,44639,51262,55732,59057,61693,63872,0),
        (34148,44642,51263,55733,59058,61693,63873,0),
        (34152,44644,51265,55734,59058,61694,63873,0),
        (34154,44646,51266,55735,59059,61694,63874,0),
        (34157,44647,51267,55736,59060,61695,63874,0),
        (34161,44650,51269,55737,59061,61695,63874,0),
        (34164,44652,51270,55738,59061,61696,63875,0),
        (34166,44654,51271,55739,59062,61697,63875,0),
        (34169,44656,51272,55740,59063,61697,63876,0),
        (34173,44658,51274,55741,59063,61698,63877,0),
        (34176,44660,51275,55741,59064,61698,63877,0),
        (34178,44662,51276,55743,59065,61699,63877,0),
        (34182,44664,51278,55743,59066,61699,63878,0),
        (34185,44666,51279,55744,59066,61700,63878,0),
        (34187,44668,51280,55745,59067,61701,63879,0),
        (34190,44670,51282,55746,59068,61701,63879,0),
        (34194,44672,51283,55747,59068,61702,63880,0),
        (34197,44674,51284,55748,59069,61702,63880,0),
        (34199,44676,51286,55749,59070,61703,63881,0),
        (34203,44678,51287,55750,59071,61703,63881,0),
        (34206,44680,51288,55751,59071,61704,63882,0),
        (34208,44682,51289,55752,59072,61705,63882,0),
        (34211,44685,51291,55753,59073,61705,63883,0),
        (34215,44686,51292,55753,59073,61706,63883,0),
        (34218,44688,51293,55754,59074,61707,63884,0),
        (34220,44690,51295,55755,59075,61707,63884,0),
        (34224,44692,51296,55756,59076,61708,63885,0),
        (34227,44694,51297,55757,59076,61708,63885,0),
        (34229,44696,51298,55758,59077,61709,63886,0),
        (34232,44699,51300,55759,59078,61709,63886,0),
        (34236,44700,51301,55760,59078,61710,63887,0),
        (34239,44702,51302,55761,59079,61711,63887,0),
        (34241,44704,51304,55762,59080,61711,63888,0),
        (34245,44707,51305,55763,59081,61712,63888,0),
        (34248,44708,51306,55764,59081,61712,63889,0),
        (34250,44710,51307,55765,59082,61713,63889,0),
        (34253,44713,51309,55766,59083,61713,63890,0),
        (34257,44715,51310,55766,59083,61714,63890,0),
        (34260,44716,51311,55767,59084,61715,63891,0),
        (34262,44718,51313,55768,59085,61715,63891,0),
        (34266,44721,51314,55769,59086,61716,63892,0),
        (34269,44722,51315,55770,59086,61716,63892,0),
        (34271,44724,51316,55771,59087,61717,63893,0),
        (34274,44727,51318,55772,59088,61717,63893,0),
        (34278,44729,51319,55773,59088,61718,63894,0),
        (34281,44730,51320,55774,59089,61719,63894,0),
        (34283,44732,51322,55775,59090,61719,63895,0),
        (34287,44735,51323,55776,59091,61720,63895,0),
        (34290,44737,51324,55777,59091,61720,63896,0),
        (34293,44738,51325,55778,59092,61721,63896,0),
        (34295,44741,51327,55779,59093,61722,63896,0),
        (34299,44743,51328,55779,59093,61722,63897,0),
        (34302,44744,51329,55780,59094,61723,63897,0),
        (34304,44746,51331,55781,59095,61723,63898,0),
        (34308,44749,51332,55782,59095,61724,63898,0),
        (34311,44751,51333,55783,59096,61725,63899,0),
        (34314,44752,51334,55784,59097,61725,63899,0),
        (34316,44755,51336,55785,59098,61726,63900,0),
        (34320,44757,51337,55786,59098,61726,63900,0),
        (34323,44759,51338,55787,59099,61727,63901,0),
        (34325,44760,51340,55788,59100,61727,63901,0),
        (34329,44763,51341,55789,59100,61728,63902,0),
        (34332,44765,51342,55789,59101,61729,63902,0),
        (34335,44766,51343,55791,59102,61729,63903,0),
        (34337,44769,51345,55791,59103,61730,63903,0),
        (34341,44771,51346,55792,59103,61730,63904,0),
        (34344,44773,51347,55793,59104,61731,63904,0),
        (34346,44774,51349,55794,59105,61731,63905,0),
        (34350,44777,51350,55795,59105,61732,63905,0),
        (34353,44779,51351,55796,59106,61733,63906,0),
        (34356,44781,51352,55797,59107,61733,63906,0),
        (34358,44783,51354,55798,59108,61734,63907,0),
        (34362,44785,51355,55799,59108,61734,63907,0),
        (34365,44787,51356,55799,59109,61735,63908,0),
        (34367,44788,51358,55801,59110,61735,63908,0),
        (34371,44791,51359,55802,59110,61736,63909,0),
        (34374,44793,51360,55802,59111,61737,63909,0),
        (34377,44795,51361,55804,59112,61737,63910,0),
        (34379,44797,51363,55804,59113,61738,63910,0),
        (34383,44799,51364,55805,59113,61738,63911,0),
        (34386,44801,51365,55806,59114,61739,63911,0),
        (34388,44802,51367,55807,59115,61739,63912,0),
        (34392,44805,51368,55808,59115,61740,63912,0),
        (34395,44807,51369,55809,59116,61741,63913,0),
        (34398,44809,51370,55810,59117,61741,63913,0),
        (34400,44811,51372,55811,59118,61742,63913,0),
        (34404,44813,51373,55812,59118,61742,63914,0),
        (34407,44815,51374,55812,59119,61743,63915,0),
        (34409,44816,51376,55814,59120,61744,63915,0),
        (34413,44819,51377,55814,59120,61744,63915,0),
        (34416,44821,51378,55815,59121,61745,63916,0),
        (34419,44823,51380,55816,59122,61745,63916,0),
        (34422,44825,51381,55817,59123,61746,63917,0),
        (34425,44827,51382,55818,59123,61747,63918,0),
        (34428,44829,51383,55819,59124,61747,63918,0),
        (34430,44831,51385,55820,59125,61748,63918,0),
        (34434,44833,51386,55821,59125,61748,63919,0),
        (34437,44835,51387,55822,59126,61749,63919,0),
        (34440,44837,51389,55823,59127,61749,63920,0),
        (34443,44839,51390,55824,59128,61750,63920,0),
        (34446,44841,51391,55824,59128,61751,63921,0),
        (34449,44843,51392,55826,59129,61751,63921,0),
        (34451,44845,51394,55826,59130,61752,63922,0),
        (34455,44847,51395,55827,59130,61752,63922,0),
        (34458,44849,51396,55828,59131,61753,63923,0),
        (34461,44851,51398,55829,59132,61753,63923,0),
        (34464,44853,51399,55830,59133,61754,63924,0),
        (34467,44855,51400,55831,59133,61755,63924,0),
        (34470,44857,51401,55832,59134,61755,63925,0),
        (34472,44859,51403,55833,59135,61756,63925,0),
        (34476,44861,51404,55834,59135,61756,63926,0),
        (34479,44863,51405,55835,59136,61757,63926,0),
        (34482,44865,51407,55836,59137,61757,63927,0),
        (34485,44867,51408,55837,59138,61758,63927,0),
        (34488,44869,51409,55837,59138,61759,63928,0),
        (34491,44871,51410,55839,59139,61759,63928,0),
        (34493,44873,51412,55839,59140,61760,63929,0),
        (34497,44875,51413,55840,59140,61760,63929,0),
        (34500,44877,51414,55841,59141,61761,63930,0),
        (34502,44879,51416,55842,59142,61762,63930,0),
        (34506,44881,51417,55843,59143,61762,63931,0),
        (34509,44883,51418,55844,59143,61763,63931,0),
        (34512,44885,51419,55845,59144,61763,63932,0),
        (34514,44887,51421,55846,59145,61764,63932,0),
        (34518,44889,51422,55847,59145,61764,63933,0),
        (34521,44891,51423,55847,59146,61765,63933,0),
        (34523,44892,51425,55849,59147,61766,63933,0),
        (34527,44895,51426,55849,59147,61766,63934,0),
        (34530,44897,51427,55850,59148,61767,63935,0),
        (34533,44899,51428,55851,59149,61767,63935,0),
        (34535,44901,51430,55852,59150,61768,63935,0),
        (34539,44903,51431,55853,59150,61768,63936,0),
        (34542,44905,51432,55854,59151,61769,63936,0),
        (34544,44906,51433,55855,59152,61770,63937,0),
        (34548,44909,51435,55856,59152,61770,63937,0),
        (34551,44911,51436,55857,59153,61771,63938,0),
        (34554,44913,51437,55858,59154,61771,63938,0),
        (34556,44915,51439,55859,59155,61772,63939,0),
        (34560,44917,51440,55859,59155,61772,63939,0),
        (34563,44919,51441,55860,59156,61773,63940,0),
        (34565,44920,51442,55861,59157,61774,63940,0),
        (34569,44923,51444,55862,59157,61774,63941,0),
        (34572,44925,51445,55863,59158,61775,63941,0),
        (34575,44926,51446,55864,59159,61775,63942,0),
        (34577,44929,51447,55865,59160,61776,63942,0),
        (34581,44931,51449,55866,59160,61776,63943,0),
        (34584,44933,51450,55867,59161,61777,63943,0),
        (34586,44934,51451,55868,59162,61778,63944,0),
        (34590,44937,51452,55869,59162,61778,63944,0),
        (34593,44939,51454,55869,59163,61779,63945,0),
        (34596,44940,51455,55871,59164,61779,63945,0),
        (34598,44943,51456,55871,59165,61780,63946,0),
        (34602,44945,51458,55872,59165,61780,63946,0),
        (34605,44946,51459,55873,59166,61781,63947,0),
        (34607,44948,51460,55874,59167,61782,63947,0),
        (34611,44951,51461,55875,59167,61782,63948,0),
        (34614,44953,51463,55876,59168,61783,63948,0),
        (34616,44954,51464,55877,59169,61783,63949,0),
        (34619,44957,51465,55878,59170,61784,63949,0),
        (34623,44959,51466,55879,59170,61784,63950,0),
        (34626,44960,51468,55879,59171,61785,63950,0),
        (34628,44962,51469,55881,59172,61786,63950,0),
        (34632,44965,51470,55881,59172,61786,63951,0),
        (34635,44966,51471,55882,59173,61787,63952,0),
        (34637,44968,51473,55883,59174,61788,63952,0),
        (34640,44971,51474,55884,59174,61788,63952,0),
        (34644,44973,51475,55885,59175,61789,63953,0),
        (34647,44974,51476,55886,59176,61789,63953,0),
        (34649,44976,51478,55887,59177,61790,63954,0),
        (34653,44979,51479,55888,59177,61790,63954,0),
        (34656,44980,51480,55889,59178,61791,63955,0),
        (34658,44982,51482,55890,59179,61792,63955,0),
        (34661,44985,51483,55891,59179,61792,63956,0),
        (34665,44986,51484,55891,59180,61793,63956,0),
        (34667,44988,51485,55892,59181,61793,63957,0),
        (34670,44990,51487,55893,59182,61794,63957,0),
        (34674,44992,51488,55894,59182,61794,63958,0),
        (34677,44994,51489,55895,59183,61795,63958,0),
        (34679,44996,51490,55896,59184,61796,63959,0),
        (34682,44999,51492,55897,59184,61796,63959,0),
        (34686,45000,51493,55898,59185,61797,63960,0),
        (34688,45002,51494,55899,59186,61797,63960,0),
        (34691,45004,51496,55900,59187,61798,63961,0),
        (34695,45006,51497,55901,59187,61798,63961,0),
        (34698,45008,51498,55901,59188,61799,63962,0),
        (34700,45010,51499,55903,59189,61800,63962,0),
        (34703,45012,51501,55903,59189,61800,63963,0),
        (34707,45014,51502,55904,59190,61801,63963,0),
        (34709,45016,51503,55905,59191,61801,63964,0),
        (34712,45018,51505,55906,59192,61802,63964,0),
        (34716,45020,51506,55907,59192,61802,63965,0),
        (34718,45022,51507,55908,59193,61803,63965,0),
        (34721,45024,51508,55909,59194,61804,63966,0),
        (34724,45026,51510,55910,59194,61804,63966,0),
        (34728,45028,51511,55911,59195,61805,63967,0),
        (34730,45030,51512,55911,59196,61805,63967,0),
        (34733,45031,51514,55913,59196,61806,63967,0),
        (34737,45034,51515,55913,59197,61806,63968,0),
        (34739,45036,51516,55914,59198,61807,63969,0),
        (34742,45037,51517,55915,59199,61808,63969,0),
        (34745,45040,51519,55916,59199,61808,63969,0),
        (34749,45042,51520,55917,59200,61809,63970,0),
        (34751,45044,51521,55918,59201,61809,63970,0),
        (34754,45045,51523,55919,59201,61810,63971,0),
        (34758,45048,51524,55920,59202,61810,63971,0),
        (34760,45050,51525,55921,59203,61811,63972,0),
        (34763,45051,51526,55922,59204,61812,63972,0),
        (34766,45054,51528,55923,59204,61812,63973,0),
        (34769,45056,51529,55923,59205,61813,63973,0),
        (34772,45057,51530,55924,59206,61813,63974,0),
        (34775,45059,51532,55925,59206,61814,63974,0),
        (34779,45062,51533,55926,59207,61814,63975,0),
        (34781,45063,51534,55927,59208,61815,63975,0),
        (34784,45065,51535,55928,59209,61816,63976,0),
        (34786,45068,51537,55929,59209,61816,63976,0),
        (34790,45069,51538,55930,59210,61817,63977,0),
        (34793,45071,51539,55931,59211,61817,63977,0),
        (34796,45073,51540,55932,59211,61818,63978,0),
        (34800,45075,51542,55933,59212,61819,63978,0),
        (34802,45077,51543,55933,59213,61819,63979,0),
        (34805,45079,51544,55935,59213,61820,63979,0),
        (34807,45081,51545,55935,59214,61820,63980,0),
        (34811,45083,51547,55936,59215,61821,63980,0),
        (34814,45085,51548,55937,59216,61822,63981,0),
        (34816,45087,51549,55938,59216,61822,63981,0),
        (34820,45089,51550,55939,59217,61823,63981,0),
        (34823,45091,51552,55940,59217,61823,63982,0),
        (34826,45093,51553,55941,59218,61824,63983,0),
        (34828,45095,51554,55942,59219,61824,63983,0),
        (34832,45097,51555,55943,59220,61825,63984,0),
        (34835,45099,51557,55943,59221,61826,63984,0),
        (34837,45100,51558,55945,59221,61826,63984,0),
        (34841,45103,51559,55945,59222,61827,63985,0),
        (34844,45105,51560,55946,59222,61827,63985,0),
        (34847,45106,51562,55947,59223,61828,63986,0),
        (34849,45109,51563,55948,59224,61828,63986,0),
        (34853,45111,51564,55949,59225,61829,63987,0),
        (34856,45112,51565,55950,59226,61830,63987,0),
        (34858,45114,51567,55951,59226,61830,63988,0),
        (34862,45117,51568,55952,59227,61831,63988,0),
        (34865,45119,51569,55953,59227,61831,63989,0),
        (34867,45120,51570,55954,59228,61832,63989,0),
        (34870,45123,51572,55955,59229,61832,63990,0),
        (34874,45125,51573,55955,59230,61833,63990,0),
        (34877,45126,51574,55956,59230,61834,63991,0),
        (34879,45128,51576,55957,59231,61834,63991,0),
        (34883,45131,51577,55958,59232,61835,63992,0),
        (34886,45132,51578,55959,59232,61835,63992,0),
        (34888,45134,51579,55960,59233,61836,63993,0),
        (34891,45137,51581,55961,59234,61836,63993,0),
        (34895,45138,51582,55962,59234,61837,63994,0),
        (34897,45140,51583,55962,59235,61838,63994,0),
        (34900,45142,51585,55964,59236,61838,63995,0),
        (34904,45144,51586,55964,59237,61839,63995,0),
        (34907,45146,51587,55965,59237,61839,63996,0),
        (34909,45148,51588,55966,59238,61840,63996,0),
        (34912,45150,51590,55967,59239,61840,63997,0),
        (34916,45152,51591,55968,59239,61841,63997,0),
        (34918,45154,51592,55969,59240,61842,63998,0),
        (34921,45155,51594,55970,59241,61842,63998,0),
        (34925,45158,51595,55971,59242,61843,63998,0),
        (34927,45160,51596,55972,59242,61843,63999,0),
        (34930,45161,51597,55973,59243,61844,63999,0),
        (34933,45164,51599,55974,59244,61844,64000,0),
        (34937,45166,51600,55974,59244,61845,64001,0),
        (34939,45167,51601,55975,59245,61846,64001,0),
        (34942,45169,51603,55976,59246,61846,64001,0),
        (34946,45172,51604,55977,59246,61847,64002,0),
        (34948,45173,51605,55978,59247,61847,64002,0),
        (34951,45175,51606,55979,59248,61848,64003,0),
        (34953,45178,51607,55980,59249,61848,64003,0),
        (34957,45179,51609,55981,59249,61849,64004,0),
        (34960,45181,51610,55982,59250,61850,64004,0),
        (34963,45183,51611,55983,59251,61850,64005,0),
        (34967,45185,51612,55984,59251,61851,64005,0),
        (34969,45187,51614,55984,59252,61851,64006,0),
        (34972,45189,51615,55986,59253,61852,64006,0),
        (34974,45191,51616,55986,59254,61852,64007,0),
        (34978,45193,51617,55987,59254,61853,64007,0),
        (34981,45195,51619,55988,59255,61854,64008,0),
        (34983,45197,51620,55989,59256,61854,64008,0),
        (34987,45199,51621,55990,59256,61855,64009,0),
        (34990,45201,51622,55991,59257,61855,64009,0),
        (34993,45203,51624,55992,59258,61856,64010,0),
        (34995,45205,51625,55993,59259,61856,64010,0),
        (34999,45207,51626,55993,59259,61857,64011,0),
        (35002,45209,51627,55994,59260,61858,64011,0),
        (35004,45210,51629,55995,59261,61858,64012,0),
        (35008,45213,51630,55996,59261,61859,64012,0),
        (35011,45215,51631,55997,59262,61859,64013,0),
        (35013,45216,51632,55998,59263,61860,64013,0),
        (35016,45219,51634,55999,59263,61860,64013,0),
        (35020,45221,51635,56000,59264,61861,64014,0),
        (35023,45222,51636,56001,59265,61862,64014,0),
        (35025,45224,51638,56002,59266,61862,64015,0),
        (35029,45227,51639,56003,59266,61863,64015,0),
        (35032,45228,51640,56003,59267,61863,64016,0),
        (35034,45230,51641,56005,59268,61864,64016,0),
        (35037,45232,51643,56005,59268,61864,64017,0),
        (35041,45234,51644,56006,59269,61865,64017,0),
        (35043,45236,51645,56007,59270,61866,64018,0),
        (35046,45238,51647,56008,59271,61866,64018,0),
        (35050,45240,51648,56009,59271,61867,64019,0),
        (35052,45242,51649,56010,59272,61867,64019,0),
        (35055,45244,51650,56011,59273,61868,64020,0),
        (35058,45246,51652,56012,59273,61868,64020,0),
        (35062,45248,51653,56013,59274,61869,64021,0),
        (35064,45250,51654,56013,59275,61870,64021,0),
        (35067,45251,51655,56014,59275,61870,64022,0),
        (35071,45254,51657,56015,59276,61871,64022,0),
        (35073,45256,51658,56016,59277,61871,64023,0),
        (35076,45257,51659,56017,59278,61872,64023,0),
        (35078,45260,51660,56018,59278,61872,64024,0),
        (35082,45262,51662,56019,59279,61873,64024,0),
        (35085,45263,51663,56020,59280,61874,64025,0),
        (35088,45265,51664,56021,59280,61874,64025,0),
        (35091,45267,51665,56022,59281,61875,64025,0),
        (35094,45269,51666,56022,59282,61875,64026,0),
        (35097,45271,51668,56024,59282,61876,64027,0),
        (35099,45273,51669,56024,59283,61876,64027,0),
        (35103,45275,51670,56025,59284,61877,64028,0),
        (35106,45277,51671,56026,59285,61878,64028,0),
        (35108,45279,51673,56027,59285,61878,64028,0),
        (35112,45281,51674,56028,59286,61879,64029,0),
        (35115,45283,51675,56029,59286,61880,64029,0),
        (35118,45285,51676,56030,59287,61880,64030,0),
        (35120,45287,51678,56031,59288,61881,64030,0),
        (35124,45289,51679,56032,59289,61881,64031,0),
        (35127,45290,51680,56032,59290,61882,64031,0),
        (35129,45292,51682,56033,59290,61882,64032,0),
        (35133,45295,51683,56034,59291,61883,64032,0),
        (35136,45296,51684,56035,59291,61884,64033,0),
        (35138,45298,51685,56036,59292,61884,64033,0),
        (35141,45301,51687,56037,59293,61885,64034,0),
        (35145,45302,51688,56038,59294,61885,64034,0),
        (35147,45304,51689,56039,59294,61886,64035,0),
        (35150,45306,51691,56040,59295,61886,64035,0),
        (35154,45308,51692,56041,59296,61887,64036,0),
        (35156,45310,51693,56041,59296,61888,64036,0),
        (35159,45312,51694,56043,59297,61888,64037,0),
        (35162,45314,51696,56043,59298,61889,64037,0),
        (35166,45316,51697,56044,59298,61889,64038,0),
        (35168,45318,51698,56045,59299,61890,64038,0),
        (35171,45319,51699,56046,59300,61890,64039,0),
        (35175,45322,51701,56047,59301,61891,64039,0),
        (35177,45324,51702,56048,59301,61892,64040,0),
        (35180,45325,51703,56049,59302,61892,64040,0),
        (35182,45328,51704,56050,59303,61893,64040,0),
        (35186,45330,51705,56051,59303,61893,64041,0),
        (35189,45331,51707,56051,59304,61894,64042,0),
        (35192,45333,51708,56052,59305,61894,64042,0),
        (35195,45336,51709,56053,59306,61895,64042,0),
        (35198,45337,51710,56054,59306,61896,64043,0),
        (35201,45339,51712,56055,59307,61896,64043,0),
        (35203,45341,51713,56056,59308,61897,64044,0),
        (35207,45343,51714,56057,59308,61897,64044,0),
        (35210,45345,51715,56058,59309,61898,64045,0),
        (35212,45347,51717,56059,59310,61898,64045,0),
        (35216,45349,51718,56060,59310,61899,64046,0),
        (35219,45351,51719,56060,59311,61900,64046,0),
        (35221,45352,51720,56062,59312,61900,64047,0),
        (35224,45355,51722,56062,59313,61901,64047,0),
        (35228,45357,51723,56063,59313,61901,64048,0),
        (35231,45358,51724,56064,59314,61902,64048,0),
        (35233,45361,51726,56065,59315,61902,64049,0),
        (35237,45363,51727,56066,59315,61903,64049,0),
        (35240,45364,51728,56067,59316,61904,64050,0),
        (35242,45366,51730,56068,59317,61904,64050,0),
        (35246,45369,51731,56069,59317,61905,64051,0),
        (35249,45370,51732,56069,59318,61905,64051,0),
        (35251,45372,51733,56071,59319,61906,64052,0),
        (35254,45374,51735,56071,59320,61906,64052,0),
        (35258,45376,51736,56072,59320,61907,64053,0),
        (35260,45378,51737,56073,59321,61908,64053,0),
        (35263,45380,51738,56074,59322,61908,64054,0),
        (35267,45382,51739,56075,59322,61909,64054,0),
        (35269,45384,51741,56076,59323,61909,64055,0),
        (35272,45385,51742,56077,59324,61910,64055,0),
        (35275,45388,51743,56078,59325,61910,64055,0),
        (35279,45390,51744,56079,59325,61911,64056,0),
        (35281,45391,51745,56079,59326,61912,64056,0),
        (35284,45393,51747,56081,59327,61912,64057,0),
        (35288,45396,51748,56081,59327,61913,64057,0),
        (35290,45397,51749,56082,59328,61913,64058,0),
        (35293,45399,51750,56083,59329,61914,64058,0),
        (35295,45402,51752,56084,59329,61914,64059,0),
        (35299,45403,51753,56085,59330,61915,64059,0),
        (35302,45405,51754,56086,59331,61916,64060,0),
        (35304,45407,51756,56087,59332,61916,64060,0),
        (35308,45409,51757,56088,59332,61917,64061,0),
        (35311,45411,51758,56088,59333,61917,64061,0),
        (35314,45413,51759,56090,59334,61918,64062,0),
        (35316,45415,51761,56090,59334,61918,64062,0),
        (35320,45417,51762,56091,59335,61919,64063,0),
        (35323,45418,51763,56092,59336,61920,64063,0),
        (35325,45420,51765,56093,59336,61920,64064,0),
        (35329,45423,51766,56094,59337,61921,64064,0),
        (35332,45424,51767,56095,59338,61921,64065,0),
        (35334,45426,51768,56096,59339,61922,64065,0),
        (35337,45429,51769,56097,59339,61922,64066,0),
        (35341,45430,51771,56097,59340,61923,64066,0),
        (35343,45432,51772,56098,59341,61923,64067,0),
        (35346,45434,51773,56099,59341,61924,64067,0),
        (35350,45436,51774,56100,59342,61924,64067,0),
        (35352,45438,51775,56101,59343,61925,64068,0),
        (35355,45440,51777,56102,59344,61926,64068,0),
        (35358,45442,51778,56103,59344,61926,64069,0),
        (35361,45444,51779,56104,59345,61927,64070,0),
        (35364,45445,51780,56105,59346,61927,64070,0),
        (35367,45447,51782,56106,59346,61928,64070,0),
        (35371,45450,51783,56107,59347,61928,64071,0),
        (35373,45451,51784,56107,59347,61929,64071,0),
        (35376,45453,51785,56108,59348,61930,64072,0),
        (35378,45456,51787,56109,59349,61930,64072,0),
        (35382,45457,51788,56110,59350,61931,64073,0),
        (35385,45459,51789,56111,59351,61931,64073,0),
        (35387,45461,51791,56112,59351,61932,64074,0),
        (35391,45463,51792,56113,59352,61932,64074,0),
        (35394,45465,51793,56114,59352,61933,64075,0),
        (35396,45467,51794,56115,59353,61934,64075,0),
        (35399,45469,51796,56116,59354,61934,64076,0),
        (35403,45471,51797,56116,59355,61935,64076,0),
        (35406,45472,51798,56117,59355,61935,64077,0),
        (35408,45474,51799,56118,59356,61936,64077,0),
        (35412,45477,51801,56119,59357,61936,64078,0),
        (35415,45478,51802,56120,59357,61937,64078,0),
        (35417,45480,51803,56121,59358,61938,64079,0),
        (35420,45482,51804,56122,59359,61938,64079,0),
        (35424,45484,51805,56123,59359,61939,64080,0),
        (35426,45486,51807,56123,59360,61939,64080,0),
        (35429,45488,51808,56125,59361,61940,64080,0),
        (35433,45490,51809,56125,59362,61940,64081,0),
        (35435,45492,51810,56126,59362,61941,64082,0),
        (35438,45493,51811,56127,59363,61942,64082,0),
        (35440,45496,51813,56128,59364,61942,64082,0),
        (35444,45498,51814,56129,59364,61943,64083,0),
        (35447,45499,51815,56130,59365,61943,64083,0),
        (35449,45501,51817,56131,59366,61944,64084,0),
        (35453,45503,51818,56132,59366,61944,64084,0),
        (35456,45505,51819,56132,59367,61945,64085,0),
        (35459,45507,51820,56134,59368,61946,64085,0),
        (35461,45509,51822,56134,59369,61946,64086,0),
        (35465,45511,51823,56135,59369,61947,64086,0),
        (35468,45513,51824,56136,59370,61947,64087,0),
        (35470,45514,51826,56137,59371,61948,64087,0),
        (35474,45517,51827,56138,59371,61948,64088,0),
        (35477,45519,51828,56139,59372,61949,64088,0),
        (35479,45520,51829,56140,59373,61950,64089,0),
        (35482,45523,51831,56141,59373,61950,64089,0),
        (35486,45524,51832,56141,59374,61951,64090,0),
        (35488,45526,51833,56142,59375,61951,64090,0),
        (35491,45528,51834,56143,59376,61952,64091,0),
        (35495,45530,51835,56144,59376,61952,64091,0),
        (35497,45532,51836,56145,59377,61953,64092,0),
        (35500,45534,51838,56146,59378,61954,64092,0),
        (35502,45536,51839,56147,59378,61954,64092,0),
        (35506,45538,51840,56148,59379,61955,64093,0),
        (35509,45540,51841,56149,59380,61955,64093,0),
        (35512,45541,51843,56150,59380,61956,64094,0),
        (35515,45544,51844,56151,59381,61956,64094,0),
        (35518,45545,51845,56151,59382,61957,64095,0),
        (35521,45547,51846,56152,59383,61958,64095,0),
        (35523,45550,51848,56153,59383,61958,64096,0),
        (35527,45551,51849,56154,59384,61959,64096,0),
        (35530,45553,51850,56155,59385,61959,64097,0),
        (35532,45555,51852,56156,59385,61960,64097,0),
        (35536,45557,51853,56157,59386,61960,64098,0),
        (35539,45559,51854,56158,59387,61961,64098,0),
        (35541,45560,51855,56159,59387,61962,64099,0),
        (35544,45563,51857,56160,59388,61962,64099,0),
        (35548,45565,51858,56160,59389,61963,64100,0),
        (35550,45566,51859,56161,59390,61963,64100,0),
        (35553,45568,51860,56162,59390,61964,64101,0),
        (35557,45571,51861,56163,59391,61964,64101,0),
        (35559,45572,51863,56164,59391,61965,64102,0),
        (35562,45574,51864,56165,59392,61966,64102,0),
        (35564,45576,51865,56166,59393,61966,64103,0),
        (35568,45578,51866,56167,59394,61967,64103,0),
        (35571,45580,51867,56167,59394,61967,64104,0),
        (35574,45581,51869,56169,59395,61968,64104,0),
        (35577,45584,51870,56169,59396,61968,64104,0),
        (35580,45586,51871,56170,59396,61969,64105,0),
        (35583,45587,51872,56171,59397,61970,64105,0),
        (35585,45590,51874,56172,59398,61970,64106,0),
        (35589,45591,51875,56173,59398,61971,64106,0),
        (35592,45593,51876,56174,59399,61971,64107,0),
        (35594,45595,51878,56175,59400,61972,64107,0),
        (35598,45597,51879,56176,59401,61972,64108,0),
        (35601,45599,51880,56176,59401,61973,64108,0),
        (35603,45601,51881,56178,59402,61974,64109,0),
        (35606,45603,51883,56178,59403,61974,64109,0),
        (35610,45605,51884,56179,59403,61975,64110,0),
        (35612,45606,51885,56180,59404,61975,64110,0),
        (35615,45608,51886,56181,59405,61976,64111,0),
        (35619,45611,51887,56182,59405,61976,64111,0),
        (35621,45612,51889,56183,59406,61977,64112,0),
        (35624,45614,51890,56184,59407,61978,64112,0),
        (35626,45616,51891,56185,59408,61978,64113,0),
        (35630,45618,51892,56185,59408,61979,64113,0),
        (35633,45620,51893,56186,59409,61979,64114,0),
        (35635,45621,51895,56187,59410,61980,64114,0),
        (35639,45624,51896,56188,59410,61980,64114,0),
        (35642,45626,51897,56189,59411,61981,64115,0),
        (35644,45627,51898,56190,59412,61982,64116,0),
        (35647,45630,51900,56191,59412,61982,64116,0),
        (35651,45631,51901,56192,59413,61983,64117,0),
        (35653,45633,51902,56192,59414,61983,64117,0),
        (35656,45635,51904,56194,59415,61984,64117,0),
        (35660,45637,51905,56194,59415,61984,64118,0),
        (35662,45639,51906,56195,59416,61985,64118,0),
        (35665,45641,51907,56196,59417,61985,64119,0),
        (35668,45643,51909,56197,59417,61986,64119,0),
        (35672,45645,51910,56198,59418,61986,64120,0),
        (35674,45646,51911,56199,59419,61987,64120,0),
        (35677,45648,51912,56200,59419,61988,64121,0),
        (35681,45651,51913,56201,59420,61988,64121,0),
        (35683,45652,51914,56201,59421,61989,64122,0),
        (35686,45654,51916,56203,59422,61989,64122,0),
        (35688,45656,51917,56203,59422,61990,64123,0),
        (35692,45658,51918,56204,59423,61990,64123,0),
        (35695,45660,51919,56205,59424,61991,64124,0),
        (35697,45661,51921,56206,59424,61992,64124,0),
        (35701,45664,51922,56207,59425,61992,64125,0),
        (35704,45666,51923,56208,59426,61993,64125,0),
        (35706,45667,51924,56209,59426,61993,64126,0),
        (35709,45670,51926,56210,59427,61994,64126,0),
        (35713,45671,51927,56210,59428,61994,64127,0),
        (35715,45673,51928,56211,59429,61995,64127,0),
        (35718,45675,51930,56212,59429,61996,64127,0),
        (35722,45677,51931,56213,59430,61996,64128,0),
        (35724,45679,51932,56214,59430,61997,64129,0),
        (35727,45681,51933,56215,59431,61997,64129,0),
        (35729,45683,51934,56216,59432,61998,64129,0),
        (35733,45685,51936,56217,59433,61998,64130,0),
        (35736,45686,51937,56217,59433,61999,64130,0),
        (35738,45688,51938,56219,59434,62000,64131,0),
        (35742,45691,51939,56219,59435,62000,64131,0),
        (35745,45692,51940,56220,59435,62001,64132,0),
        (35747,45694,51941,56221,59436,62001,64132,0),
        (35750,45696,51943,56222,59437,62002,64133,0),
        (35754,45698,51944,56223,59437,62002,64133,0),
        (35756,45700,51945,56224,59438,62003,64134,0),
        (35759,45701,51947,56225,59439,62004,64134,0),
        (35763,45704,51948,56226,59440,62004,64135,0),
        (35765,45705,51949,56226,59440,62005,64135,0),
        (35768,45707,51950,56228,59441,62005,64136,0),
        (35771,45710,51952,56228,59442,62006,64136,0),
        (35774,45711,51953,56229,59442,62006,64137,0),
        (35777,45713,51954,56230,59443,62007,64137,0),
        (35780,45715,51955,56231,59444,62008,64138,0),
        (35783,45717,51957,56232,59444,62008,64138,0),
        (35786,45719,51958,56233,59445,62009,64139,0),
        (35789,45720,51959,56234,59446,62009,64139,0),
        (35791,45723,51960,56235,59446,62010,64139,0),
        (35795,45725,51961,56235,59447,62010,64140,0),
        (35798,45726,51962,56236,59448,62011,64140,0),
        (35800,45728,51964,56237,59449,62012,64141,0),
        (35804,45730,51965,56238,59449,62012,64141,0),
        (35807,45732,51966,56239,59450,62013,64142,0),
        (35809,45734,51967,56240,59451,62013,64142,0),
        (35812,45736,51969,56241,59451,62014,64143,0),
        (35816,45738,51970,56242,59452,62014,64143,0),
        (35818,45739,51971,56242,59453,62015,64144,0),
        (35821,45741,51973,56244,59453,62015,64144,0),
        (35825,45744,51974,56244,59454,62016,64145,0),
        (35827,45745,51975,56245,59455,62017,64145,0),
        (35830,45747,51976,56246,59456,62017,64146,0),
        (35832,45749,51978,56247,59456,62018,64146,0),
        (35836,45751,51979,56248,59457,62018,64147,0),
        (35839,45753,51980,56249,59458,62019,64147,0),
        (35841,45754,51981,56250,59458,62019,64148,0),
        (35845,45757,51982,56251,59459,62020,64148,0),
        (35848,45758,51983,56251,59460,62021,64149,0),
        (35850,45760,51985,56252,59460,62021,64149,0),
        (35853,45763,51986,56253,59461,62022,64149,0),
        (35857,45764,51987,56254,59462,62022,64150,0),
        (35859,45766,51988,56255,59463,62023,64150,0),
        (35862,45768,51990,56256,59463,62023,64151,0),
        (35866,45770,51991,56257,59464,62024,64151,0),
        (35868,45772,51992,56258,59464,62025,64152,0),
        (35871,45773,51993,56259,59465,62025,64152,0),
        (35873,45776,51995,56259,59466,62026,64153,0),
        (35877,45777,51996,56260,59466,62026,64153,0),
        (35880,45779,51997,56261,59467,62027,64154,0),
        (35882,45781,51998,56262,59468,62027,64154,0),
        (35886,45783,52000,56263,59469,62028,64155,0),
        (35889,45785,52001,56264,59469,62029,64155,0),
        (35891,45786,52002,56265,59470,62029,64156,0),
        (35894,45789,52003,56266,59471,62030,64156,0),
        (35898,45791,52004,56266,59471,62030,64157,0),
        (35900,45792,52005,56267,59472,62031,64157,0),
        (35903,45794,52007,56268,59473,62031,64158,0),
        (35907,45796,52008,56269,59473,62032,64158,0),
        (35909,45798,52009,56270,59474,62033,64159,0),
        (35912,45800,52010,56271,59475,62033,64159,0),
        (35914,45802,52012,56272,59476,62034,64159,0),
        (35918,45804,52013,56273,59476,62034,64160,0),
        (35921,45805,52014,56273,59477,62035,64161,0),
        (35923,45807,52016,56275,59478,62035,64161,0),
        (35927,45810,52017,56275,59478,62036,64161,0),
        (35930,45811,52018,56276,59479,62037,64162,0),
        (35932,45813,52019,56277,59480,62037,64162,0),
        (35935,45815,52020,56278,59480,62038,64163,0),
        (35939,45817,52022,56279,59481,62038,64163,0),
        (35941,45819,52023,56280,59482,62039,64164,0),
        (35944,45820,52024,56281,59483,62039,64164,0),
        (35948,45823,52025,56282,59483,62040,64165,0),
        (35950,45824,52026,56282,59484,62040,64165,0),
        (35953,45826,52027,56284,59485,62041,64166,0),
        (35955,45829,52029,56284,59485,62041,64166,0),
        (35959,45830,52030,56285,59486,62042,64167,0),
        (35962,45832,52031,56286,59487,62043,64167,0),
        (35964,45833,52033,56287,59487,62043,64168,0),
        (35968,45836,52034,56288,59488,62044,64168,0),
        (35971,45838,52035,56289,59489,62044,64169,0),
        (35973,45839,52036,56290,59489,62045,64169,0),
        (35976,45842,52038,56291,59490,62045,64169,0),
        (35980,45843,52039,56291,59491,62046,64170,0),
        (35982,45845,52040,56292,59492,62047,64171,0),
        (35985,45847,52041,56293,59492,62047,64171,0),
        (35989,45849,52042,56294,59493,62048,64171,0),
        (35991,45851,52043,56295,59493,62048,64172,0),
        (35994,45852,52045,56296,59494,62049,64172,0),
        (35996,45855,52046,56297,59495,62049,64173,0),
        (36000,45856,52047,56298,59496,62050,64173,0),
        (36003,45858,52048,56298,59496,62051,64174,0),
        (36005,45860,52050,56299,59497,62051,64174,0),
        (36009,45862,52051,56300,59498,62052,64175,0),
        (36012,45864,52052,56301,59498,62052,64175,0),
        (36014,45865,52053,56302,59499,62053,64176,0),
        (36017,45868,52055,56303,59500,62053,64176,0),
        (36021,45870,52056,56304,59500,62054,64177,0),
        (36023,45871,52057,56305,59501,62055,64177,0),
        (36026,45873,52058,56306,59502,62055,64178,0),
        (36030,45875,52060,56306,59502,62056,64178,0),
        (36032,45877,52061,56307,59503,62056,64179,0),
        (36035,45879,52062,56308,59504,62057,64179,0),
        (36039,45881,52063,56309,59505,62057,64180,0),
        (36041,45883,52064,56310,59505,62058,64180,0),
        (36044,45884,52065,56311,59506,62059,64181,0),
        (36046,45887,52067,56312,59507,62059,64181,0),
        (36050,45888,52068,56313,59507,62060,64182,0),
        (36053,45890,52069,56313,59508,62060,64182,0),
        (36055,45892,52071,56315,59509,62061,64182,0),
        (36059,45894,52072,56315,59509,62061,64183,0),
        (36062,45896,52073,56316,59510,62062,64183,0),
        (36064,45897,52074,56317,59511,62062,64184,0),
        (36067,45900,52076,56318,59512,62063,64184,0),
        (36071,45902,52077,56319,59512,62063,64185,0),
        (36073,45903,52078,56320,59513,62064,64185,0),
        (36076,45905,52079,56321,59514,62065,64186,0),
        (36080,45907,52080,56322,59514,62065,64186,0),
        (36082,45909,52081,56322,59515,62066,64187,0),
        (36085,45911,52082,56323,59516,62066,64187,0),
        (36087,45913,52084,56324,59516,62067,64188,0),
        (36091,45915,52085,56325,59517,62067,64188,0),
        (36094,45916,52086,56326,59518,62068,64189,0),
        (36096,45918,52088,56327,59518,62069,64189,0),
        (36100,45920,52089,56328,59519,62069,64190,0),
        (36103,45922,52090,56329,59520,62070,64190,0),
        (36105,45924,52091,56330,59521,62070,64191,0),
        (36108,45926,52093,56330,59521,62071,64191,0),
        (36111,45928,52094,56331,59522,62071,64192,0),
        (36114,45929,52095,56332,59523,62072,64192,0),
        (36117,45931,52096,56333,59523,62073,64192,0),
        (36120,45933,52097,56334,59524,62073,64193,0),
        (36123,45935,52098,56335,59525,62074,64193,0),
        (36125,45937,52100,56336,59525,62074,64194,0),
        (36128,45939,52101,56337,59526,62075,64194,0),
        (36132,45941,52102,56337,59527,62075,64195,0),
        (36134,45942,52103,56338,59528,62076,64195,0),
        (36137,45944,52105,56339,59528,62077,64196,0),
        (36141,45947,52106,56340,59529,62077,64196,0),
        (36143,45948,52107,56341,59529,62078,64197,0),
        (36146,45950,52108,56342,59530,62078,64197,0),
        (36148,45952,52110,56343,59531,62079,64198,0),
        (36152,45954,52111,56344,59531,62079,64198,0),
        (36155,45956,52112,56344,59532,62080,64199,0),
        (36157,45957,52113,56346,59533,62080,64199,0),
        (36161,45960,52114,56346,59534,62081,64200,0),
        (36164,45961,52116,56347,59534,62082,64200,0),
        (36166,45963,52117,56348,59535,62082,64201,0),
        (36169,45965,52118,56349,59536,62083,64201,0),
        (36173,45967,52119,56350,59536,62083,64202,0),
        (36175,45969,52120,56351,59537,62084,64202,0),
        (36178,45970,52122,56352,59538,62084,64202,0),
        (36182,45973,52123,56352,59538,62085,64203,0),
        (36184,45974,52124,56353,59539,62086,64203,0),
        (36187,45976,52125,56354,59540,62086,64204,0),
        (36189,45978,52127,56355,59541,62087,64204,0),
        (36193,45980,52128,56356,59541,62087,64205,0),
        (36196,45982,52129,56357,59542,62088,64205,0),
        (36198,45983,52130,56358,59543,62088,64206,0),
        (36202,45986,52131,56359,59543,62089,64206,0),
        (36205,45987,52133,56359,59544,62090,64207,0),
        (36207,45989,52134,56361,59545,62090,64207,0),
        (36210,45991,52135,56361,59545,62091,64208,0),
        (36213,45993,52136,56362,59546,62091,64208,0),
        (36216,45995,52137,56363,59547,62092,64209,0),
        (36219,45996,52139,56364,59547,62092,64209,0),
        (36222,45999,52140,56365,59548,62093,64210,0),
        (36225,46000,52141,56366,59549,62094,64210,0),
        (36228,46002,52142,56367,59550,62094,64211,0),
        (36230,46004,52144,56368,59550,62095,64211,0),
        (36234,46006,52145,56368,59551,62095,64212,0),
        (36236,46008,52146,56369,59552,62096,64212,0),
        (36239,46009,52147,56370,59552,62096,64212,0),
        (36243,46012,52148,56371,59553,62097,64213,0),
        (36245,46013,52150,56372,59553,62097,64213,0),
        (36248,46015,52151,56373,59554,62098,64214,0),
        (36250,46017,52152,56374,59555,62098,64214,0),
        (36254,46019,52153,56374,59556,62099,64215,0),
        (36257,46021,52154,56375,59556,62100,64215,0),
        (36259,46022,52156,56376,59557,62100,64216,0),
        (36263,46025,52157,56377,59558,62101,64216,0),
        (36266,46026,52158,56378,59558,62101,64217,0),
        (36268,46028,52159,56379,59559,62102,64217,0),
        (36271,46030,52161,56380,59560,62102,64218,0),
        (36275,46032,52162,56381,59560,62103,64218,0),
        (36277,46034,52163,56381,59561,62104,64219,0),
        (36280,46035,52164,56383,59562,62104,64219,0),
        (36284,46038,52165,56383,59562,62105,64219,0),
        (36286,46039,52167,56384,59563,62105,64220,0),
        (36289,46041,52168,56385,59564,62106,64221,0),
        (36291,46043,52169,56386,59565,62106,64221,0),
        (36295,46045,52170,56387,59565,62107,64222,0),
        (36298,46047,52171,56388,59566,62108,64222,0),
        (36300,46048,52173,56389,59567,62108,64222,0),
        (36304,46051,52174,56389,59567,62109,64223,0),
        (36306,46052,52175,56390,59568,62109,64223,0),
        (36309,46054,52176,56391,59569,62110,64224,0),
        (36311,46056,52178,56392,59569,62110,64224,0),
        (36315,46058,52179,56393,59570,62111,64225,0),
        (36318,46060,52180,56394,59571,62111,64225,0),
        (36320,46061,52181,56395,59571,62112,64226,0),
        (36324,46064,52182,56396,59572,62112,64226,0),
        (36327,46065,52183,56396,59573,62113,64227,0),
        (36329,46067,52185,56398,59574,62114,64227,0),
        (36332,46069,52186,56398,59574,62114,64228,0),
        (36336,46071,52187,56399,59575,62115,64228,0),
        (36338,46073,52188,56400,59576,62115,64229,0),
        (36341,46074,52190,56401,59576,62116,64229,0),
        (36345,46077,52191,56402,59577,62116,64229,0),
        (36347,46078,52192,56403,59577,62117,64230,0),
        (36350,46080,52193,56404,59578,62118,64231,0),
        (36352,46082,52195,56404,59579,62118,64231,0),
        (36356,46084,52196,56405,59580,62119,64232,0),
        (36359,46086,52197,56406,59580,62119,64232,0),
        (36361,46087,52198,56407,59581,62120,64232,0),
        (36365,46090,52199,56408,59582,62120,64233,0),
        (36367,46091,52200,56409,59582,62121,64233,0),
        (36370,46093,52201,56410,59583,62122,64234,0),
        (36372,46095,52203,56411,59584,62122,64234,0),
        (36376,46097,52204,56411,59584,62123,64235,0),
        (36379,46099,52205,56412,59585,62123,64235,0),
        (36381,46100,52207,56413,59586,62124,64236,0),
        (36385,46103,52208,56414,59586,62124,64236,0),
        (36388,46104,52209,56415,59587,62125,64237,0),
        (36390,46106,52210,56416,59588,62125,64237,0),
        (36393,46108,52212,56417,59589,62126,64238,0),
        (36397,46110,52213,56418,59589,62126,64238,0),
        (36399,46111,52214,56418,59590,62127,64239,0),
        (36402,46113,52215,56419,59591,62128,64239,0),
        (36405,46116,52216,56420,59591,62128,64239,0),
        (36408,46117,52217,56421,59592,62129,64240,0),
        (36411,46119,52218,56422,59593,62129,64240,0),
        (36413,46121,52220,56423,59593,62130,64241,0),
        (36417,46123,52221,56424,59594,62130,64242,0),
        (36419,46124,52222,56424,59595,62131,64242,0),
        (36422,46126,52224,56426,59595,62132,64242,0),
        (36426,46128,52225,56426,59596,62132,64243,0),
        (36428,46130,52226,56427,59597,62133,64243,0),
        (36431,46132,52227,56428,59598,62133,64244,0),
        (36433,46134,52228,56429,59598,62134,64244,0),
        (36437,46136,52229,56430,59599,62134,64245,0),
        (36440,46137,52231,56431,59600,62135,64245,0),
        (36442,46139,52232,56432,59600,62136,64246,0),
        (36446,46141,52233,56433,59601,62136,64246,0),
        (36449,46143,52234,56433,59601,62137,64247,0),
        (36451,46145,52235,56434,59602,62137,64247,0),
        (36454,46147,52237,56435,59603,62138,64248,0),
        (36457,46149,52238,56436,59604,62138,64248,0),
        (36460,46150,52239,56437,59604,62139,64249,0),
        (36463,46152,52241,56438,59605,62139,64249,0),
        (36466,46154,52242,56439,59606,62140,64249,0),
        (36469,46156,52243,56439,59606,62141,64250,0),
        (36471,46157,52244,56441,59607,62141,64250,0),
        (36474,46160,52245,56441,59608,62142,64251,0),
        (36478,46162,52246,56442,59608,62142,64251,0),
        (36480,46163,52247,56443,59609,62143,64252,0),
        (36483,46165,52249,56444,59610,62143,64252,0),
        (36487,46167,52250,56445,59610,62144,64253,0),
        (36489,46169,52251,56446,59611,62145,64253,0),
        (36492,46170,52252,56447,59612,62145,64254,0),
        (36494,46173,52254,56447,59613,62146,64254,0),
        (36498,46174,52255,56448,59613,62146,64255,0),
        (36501,46176,52256,56449,59614,62147,64255,0),
        (36503,46178,52257,56450,59615,62147,64256,0),
        (36507,46180,52258,56451,59615,62148,64256,0),
        (36509,46182,52260,56452,59616,62149,64257,0),
        (36512,46183,52261,56453,59617,62149,64257,0),
        (36514,46186,52262,56454,59617,62150,64257,0),
        (36518,46187,52263,56454,59618,62150,64258,0),
        (36521,46189,52264,56455,59619,62151,64259,0),
        (36523,46190,52266,56456,59619,62151,64259,0),
        (36527,46193,52267,56457,59620,62152,64259,0),
        (36530,46194,52268,56458,59621,62152,64260,0),
        (36532,46196,52269,56459,59622,62153,64260,0),
        (36535,46199,52271,56460,59622,62153,64261,0),
        (36538,46200,52272,56461,59623,62154,64261,0),
        (36541,46202,52273,56461,59624,62155,64262,0),
        (36544,46203,52274,56462,59624,62155,64262,0),
        (36547,46206,52275,56463,59625,62156,64263,0),
        (36550,46207,52276,56464,59625,62156,64263,0),
        (36552,46209,52277,56465,59626,62157,64264,0),
        (36555,46211,52279,56466,59627,62157,64264,0),
        (36559,46213,52280,56467,59628,62158,64265,0),
        (36561,46215,52281,56467,59628,62159,64265,0),
        (36564,46216,52283,56469,59629,62159,64266,0),
        (36568,46219,52284,56469,59630,62160,64266,0),
        (36570,46220,52285,56470,59630,62160,64267,0),
        (36573,46222,52286,56471,59631,62161,64267,0),
        (36575,46224,52287,56472,59632,62161,64267,0),
        (36579,46226,52288,56473,59632,62162,64268,0),
        (36581,46227,52289,56474,59633,62163,64268,0),
        (36584,46229,52291,56475,59634,62163,64269,0),
        (36588,46231,52292,56475,59634,62164,64269,0),
        (36590,46233,52293,56476,59635,62164,64270,0),
        (36593,46235,52294,56477,59636,62165,64270,0),
        (36595,46237,52296,56478,59637,62165,64271,0),
        (36599,46239,52297,56479,59637,62166,64271,0),
        (36602,46240,52298,56480,59638,62166,64272,0),
        (36604,46242,52299,56481,59639,62167,64272,0),
        (36608,46244,52301,56482,59639,62167,64273,0),
        (36610,46246,52302,56482,59640,62168,64273,0),
        (36613,46247,52303,56483,59641,62169,64274,0),
        (36616,46250,52304,56484,59641,62169,64274,0),
        (36619,46251,52305,56485,59642,62170,64275,0),
        (36622,46253,52306,56486,59643,62170,64275,0),
        (36624,46255,52308,56487,59643,62171,64275,0),
        (36628,46257,52309,56488,59644,62171,64276,0),
        (36631,46259,52310,56488,59645,62172,64277,0),
        (36633,46260,52311,56490,59645,62173,64277,0),
        (36636,46263,52313,56490,59646,62173,64277,0),
        (36640,46264,52314,56491,59647,62174,64278,0),
        (36642,46266,52315,56492,59648,62174,64278,0),
        (36645,46267,52316,56493,59648,62175,64279,0),
        (36648,46270,52317,56494,59649,62175,64279,0),
        (36651,46271,52318,56495,59649,62176,64280,0),
        (36653,46273,52319,56496,59650,62176,64280,0),
        (36656,46275,52321,56496,59651,62177,64281,0),
        (36660,46277,52322,56497,59651,62177,64281,0),
        (36662,46279,52323,56498,59652,62178,64282,0),
        (36665,46280,52325,56499,59653,62179,64282,0),
        (36669,46283,52326,56500,59654,62179,64283,0),
        (36671,46284,52327,56501,59654,62180,64283,0),
        (36674,46286,52328,56502,59655,62180,64284,0),
        (36676,46288,52329,56503,59656,62181,64284,0),
        (36680,46290,52330,56503,59656,62181,64285,0),
        (36682,46291,52331,56504,59657,62182,64285,0),
        (36685,46293,52333,56505,59658,62183,64285,0),
        (36689,46295,52334,56506,59658,62183,64286,0),
        (36691,46297,52335,56507,59659,62184,64286,0),
        (36694,46299,52336,56508,59660,62184,64287,0),
        (36696,46301,52338,56509,59660,62185,64287,0),
        (36700,46303,52339,56509,59661,62185,64288,0),
        (36703,46304,52340,56510,59662,62186,64288,0),
        (36705,46306,52341,56511,59662,62186,64289,0),
        (36709,46308,52342,56512,59663,62187,64289,0),
        (36711,46310,52343,56513,59664,62188,64290,0),
        (36714,46311,52345,56514,59665,62188,64290,0),
        (36716,46314,52346,56515,59665,62189,64291,0),
        (36720,46315,52347,56516,59666,62189,64291,0),
        (36723,46317,52348,56516,59667,62190,64292,0),
        (36725,46319,52350,56517,59667,62190,64292,0),
        (36729,46321,52351,56518,59668,62191,64292,0),
        (36732,46323,52352,56519,59668,62192,64293,0),
        (36734,46324,52353,56520,59669,62192,64293,0),
        (36737,46327,52354,56521,59670,62193,64294,0),
        (36740,46328,52356,56522,59671,62193,64295,0),
        (36743,46330,52357,56522,59671,62194,64295,0),
        (36745,46331,52358,56524,59672,62194,64295,0),
        (36749,46334,52359,56524,59673,62195,64296,0),
        (36752,46335,52360,56525,59673,62196,64296,0),
        (36754,46337,52361,56526,59674,62196,64297,0),
        (36757,46339,52363,56527,59675,62197,64297,0),
        (36760,46341,52364,56528,59675,62197,64298,0),
        (36763,46343,52365,56529,59676,62198,64298,0),
        (36765,46344,52366,56530,59677,62198,64299,0),
        (36769,46346,52368,56530,59677,62199,64299,0),
        (36772,46348,52369,56531,59678,62199,64300,0),
        (36774,46350,52370,56532,59679,62200,64300,0),
        (36777,46352,52371,56533,59679,62200,64301,0),
        (36781,46354,52372,56534,59680,62201,64301,0),
        (36783,46355,52373,56535,59681,62202,64302,0),
        (36786,46357,52375,56536,59682,62202,64302,0),
        (36789,46359,52376,56537,59682,62203,64302,0),
        (36792,46361,52377,56537,59683,62203,64303,0),
        (36794,46362,52378,56538,59684,62204,64303,0),
        (36797,46365,52380,56539,59684,62204,64304,0),
        (36801,46366,52381,56540,59685,62205,64304,0),
        (36803,46368,52382,56541,59686,62206,64305,0),
        (36806,46370,52383,56542,59686,62206,64305,0),
        (36809,46372,52384,56543,59687,62207,64306,0),
        (36812,46374,52385,56543,59688,62207,64306,0),
        (36815,46375,52386,56544,59688,62208,64307,0),
        (36817,46377,52388,56545,59689,62208,64307,0),
        (36821,46379,52389,56546,59690,62209,64308,0),
        (36823,46381,52390,56547,59691,62209,64308,0),
        (36826,46383,52392,56548,59691,62210,64309,0),
        (36830,46385,52393,56549,59692,62210,64309,0),
        (36832,46386,52394,56549,59693,62211,64310,0),
        (36835,46388,52395,56551,59693,62212,64310,0),
        (36838,46390,52396,56551,59694,62212,64310,0),
        (36841,46392,52397,56552,59694,62213,64311,0),
        (36843,46393,52398,56553,59695,62213,64311,0),
        (36846,46396,52400,56554,59696,62214,64312,0),
        (36850,46397,52401,56555,59696,62214,64312,0),
        (36852,46399,52402,56556,59697,62215,64313,0),
        (36855,46401,52404,56557,59698,62216,64313,0),
        (36858,46403,52405,56557,59699,62216,64314,0),
        (36861,46404,52406,56558,59699,62217,64314,0),
        (36863,46406,52407,56559,59700,62217,64315,0),
        (36866,46408,52408,56560,59701,62218,64315,0),
        (36870,46410,52409,56561,59701,62218,64316,0),
        (36872,46412,52410,56562,59702,62219,64316,0),
        (36875,46413,52412,56563,59703,62219,64317,0),
        (36879,46416,52413,56564,59703,62220,64317,0),
        (36881,46417,52414,56564,59704,62221,64318,0),
        (36884,46419,52415,56565,59705,62221,64318,0),
        (36886,46421,52417,56566,59705,62222,64318,0),
        (36890,46423,52418,56567,59706,62222,64319,0),
        (36892,46424,52419,56568,59707,62223,64320,0),
        (36895,46426,52420,56569,59707,62223,64320,0),
        (36899,46428,52421,56570,59708,62224,64320,0),
        (36901,46430,52422,56570,59709,62225,64321,0),
        (36904,46431,52423,56571,59710,62225,64321,0),
        (36906,46434,52425,56572,59710,62226,64322,0),
        (36910,46435,52426,56573,59711,62226,64322,0),
        (36912,46437,52427,56574,59712,62227,64323,0),
        (36915,46439,52429,56575,59712,62227,64323,0),
        (36919,46441,52430,56576,59713,62228,64324,0),
        (36921,46443,52431,56576,59713,62228,64324,0),
        (36924,46444,52432,56578,59714,62229,64325,0),
        (36926,46446,52433,56578,59715,62229,64325,0),
        (36930,46448,52434,56579,59715,62230,64326,0),
        (36932,46450,52435,56580,59716,62231,64326,0),
        (36935,46451,52437,56581,59717,62231,64327,0),
        (36939,46454,52438,56582,59718,62232,64327,0),
        (36941,46455,52439,56582,59718,62232,64328,0),
        (36944,46457,52440,56584,59719,62233,64328,0),
        (36946,46459,52442,56584,59720,62233,64328,0),
        (36950,46461,52443,56585,59720,62234,64329,0),
        (36952,46462,52444,56586,59721,62235,64329,0),
        (36955,46464,52445,56587,59722,62235,64330,0),
        (36959,46466,52446,56588,59722,62236,64330,0),
        (36961,46468,52447,56589,59723,62236,64331,0),
        (36964,46469,52448,56590,59724,62237,64331,0),
        (36966,46472,52450,56590,59724,62237,64332,0),
        (36970,46473,52451,56591,59725,62238,64332,0),
        (36972,46475,52452,56592,59726,62238,64333,0),
        (36975,46476,52453,56593,59726,62239,64333,0),
        (36979,46479,52454,56594,59727,62239,64334,0),
        (36981,46480,52456,56595,59728,62240,64334,0),
        (36984,46482,52457,56596,59729,62241,64335,0),
        (36986,46484,52458,56597,59729,62241,64335,0),
        (36990,46486,52459,56597,59730,62242,64336,0),
        (36992,46488,52460,56598,59731,62242,64336,0),
        (36995,46489,52462,56599,59731,62243,64336,0),
        (36999,46491,52463,56600,59732,62243,64337,0),
        (37001,46493,52464,56601,59732,62244,64337,0),
        (37004,46495,52465,56602,59733,62245,64338,0),
        (37006,46497,52466,56603,59734,62245,64338,0),
        (37010,46499,52467,56603,59734,62246,64339,0),
        (37012,46500,52468,56604,59735,62246,64339,0),
        (37015,46502,52470,56605,59736,62247,64340,0),
        (37019,46504,52471,56606,59737,62247,64340,0),
        (37021,46506,52472,56607,59737,62248,64341,0),
        (37024,46507,52473,56608,59738,62248,64341,0),
        (37026,46510,52475,56609,59739,62249,64342,0),
        (37030,46511,52476,56609,59739,62249,64342,0),
        (37032,46513,52477,56610,59740,62250,64343,0),
        (37035,46514,52478,56611,59741,62251,64343,0),
        (37039,46517,52479,56612,59741,62251,64343,0),
        (37041,46518,52480,56613,59742,62252,64344,0),
        (37044,46520,52481,56614,59743,62252,64344,0),
        (37046,46522,52483,56615,59743,62253,64345,0),
        (37050,46524,52484,56615,59744,62253,64345,0),
        (37052,46525,52485,56616,59745,62254,64346,0),
        (37055,46527,52487,56617,59745,62255,64346,0),
        (37059,46529,52488,56618,59746,62255,64347,0),
        (37061,46531,52489,56619,59747,62256,64347,0),
        (37064,46532,52490,56620,59748,62256,64348,0),
        (37066,46535,52491,56621,59748,62257,64348,0),
        (37070,46536,52492,56621,59749,62257,64349,0),
        (37072,46538,52493,56622,59750,62258,64349,0),
        (37075,46540,52495,56623,59750,62258,64350,0),
        (37079,46542,52496,56624,59751,62259,64350,0),
        (37081,46543,52497,56625,59751,62260,64351,0),
        (37084,46545,52498,56626,59752,62260,64351,0),
        (37086,46547,52500,56627,59753,62261,64351,0),
        (37090,46549,52501,56628,59753,62261,64352,0),
        (37092,46551,52502,56628,59754,62262,64352,0),
        (37095,46552,52503,56629,59755,62262,64353,0),
        (37099,46554,52504,56630,59756,62263,64353,0),
        (37101,46556,52505,56631,59756,62263,64354,0),
        (37104,46558,52506,56632,59757,62264,64354,0),
        (37106,46560,52508,56633,59758,62264,64355,0),
        (37110,46562,52509,56634,59758,62265,64355,0),
        (37112,46563,52510,56634,59759,62266,64356,0),
        (37115,46565,52511,56635,59760,62266,64356,0),
        (37119,46567,52512,56636,59760,62267,64357,0),
        (37121,46569,52514,56637,59761,62267,64357,0),
        (37124,46570,52515,56638,59762,62268,64358,0),
        (37126,46572,52516,56639,59762,62268,64358,0),
        (37130,46574,52517,56640,59763,62269,64359,0),
        (37132,46576,52518,56640,59764,62270,64359,0),
        (37135,46577,52520,56642,59764,62270,64359,0),
        (37138,46580,52521,56642,59765,62271,64360,0),
        (37141,46581,52522,56643,59766,62271,64360,0),
        (37143,46583,52523,56644,59766,62272,64361,0),
        (37146,46585,52524,56645,59767,62272,64361,0),
        (37150,46587,52525,56646,59768,62273,64362,0),
        (37152,46588,52526,56646,59769,62273,64362,0),
        (37155,46590,52528,56648,59769,62274,64363,0),
        (37158,46592,52529,56648,59770,62274,64363,0),
        (37161,46594,52530,56649,59770,62275,64364,0),
        (37163,46595,52531,56650,59771,62276,64364,0),
        (37166,46598,52533,56651,59772,62276,64365,0),
        (37170,46599,52534,56652,59772,62277,64365,0),
        (37172,46601,52535,56652,59773,62277,64366,0),
        (37175,46602,52536,56654,59774,62278,64366,0),
        (37178,46605,52537,56654,59774,62278,64366,0),
        (37181,46606,52538,56655,59775,62279,64367,0),
        (37183,46608,52539,56656,59776,62280,64367,0),
        (37186,46610,52541,56657,59777,62280,64368,0),
        (37189,46612,52542,56658,59777,62280,64369,0),
        (37192,46613,52543,56659,59778,62281,64369,0),
        (37194,46615,52544,56660,59779,62282,64369,0),
        (37198,46617,52546,56660,59779,62282,64370,0),
        (37201,46619,52547,56661,59780,62283,64370,0),
        (37203,46620,52548,56662,59781,62283,64371,0),
        (37206,46623,52549,56663,59781,62284,64371,0),
        (37209,46624,52550,56664,59782,62284,64372,0),
        (37212,46626,52551,56665,59783,62285,64372,0),
        (37214,46627,52553,56666,59783,62286,64373,0),
        (37218,46630,52554,56666,59784,62286,64373,0),
        (37221,46631,52555,56667,59785,62287,64374,0),
        (37223,46633,52556,56668,59785,62287,64374,0),
        (37226,46635,52557,56669,59786,62288,64374,0),
        (37229,46637,52558,56670,59787,62288,64375,0),
        (37232,46638,52559,56671,59787,62289,64375,0),
        (37234,46640,52561,56672,59788,62289,64376,0),
        (37238,46642,52562,56672,59789,62290,64376,0),
        (37240,46644,52563,56673,59789,62291,64377,0),
        (37243,46645,52564,56674,59790,62291,64377,0),
        (37245,46648,52566,56675,59791,62292,64378,0),
        (37249,46649,52567,56676,59791,62292,64378,0),
        (37252,46651,52568,56677,59792,62293,64379,0),
        (37254,46652,52569,56678,59793,62293,64379,0),
        (37258,46655,52570,56678,59793,62294,64380,0),
        (37260,46656,52571,56679,59794,62295,64380,0),
        (37263,46658,52572,56680,59795,62295,64381,0),
        (37265,46660,52574,56681,59795,62296,64381,0),
        (37269,46662,52575,56682,59796,62296,64382,0),
        (37271,46663,52576,56683,59797,62297,64382,0),
        (37274,46665,52577,56684,59798,62297,64382,0),
        (37278,46667,52578,56685,59798,62298,64383,0),
        (37280,46669,52580,56685,59799,62298,64383,0),
        (37283,46670,52581,56686,59800,62299,64384,0),
        (37285,46673,52582,56687,59800,62299,64384,0),
        (37289,46674,52583,56688,59801,62300,64385,0),
        (37291,46676,52584,56689,59802,62301,64385,0),
        (37294,46677,52586,56690,59802,62301,64386,0),
        (37298,46680,52587,56691,59803,62302,64386,0),
        (37300,46681,52588,56691,59803,62302,64387,0),
        (37302,46683,52589,56692,59804,62303,64387,0),
        (37305,46685,52590,56693,59805,62303,64388,0),
        (37309,46687,52591,56694,59805,62304,64388,0),
        (37311,46688,52592,56695,59806,62304,64389,0),
        (37314,46690,52594,56696,59807,62305,64389,0),
        (37317,46692,52595,56697,59808,62305,64389,0),
        (37320,46694,52596,56697,59808,62306,64390,0),
        (37322,46695,52597,56698,59809,62307,64390,0),
        (37325,46697,52599,56699,59810,62307,64391,0),
        (37329,46699,52600,56700,59810,62308,64391,0),
        (37331,46701,52601,56701,59811,62308,64392,0),
        (37333,46702,52602,56702,59812,62309,64392,0),
        (37337,46705,52603,56703,59812,62309,64393,0),
        (37340,46706,52604,56703,59813,62310,64393,0),
        (37342,46708,52605,56704,59814,62311,64394,0),
        (37345,46710,52607,56705,59814,62311,64394,0),
        (37348,46711,52608,56706,59815,62311,64395,0),
        (37351,46713,52609,56707,59816,62312,64395,0),
        (37353,46715,52610,56708,59816,62313,64396,0),
        (37357,46717,52611,56709,59817,62313,64396,0),
        (37359,46718,52612,56709,59818,62314,64397,0),
        (37362,46720,52613,56710,59818,62314,64397,0),
        (37364,46722,52615,56711,59819,62315,64397,0),
        (37368,46724,52616,56712,59820,62315,64398,0),
        (37371,46725,52617,56713,59821,62316,64398,0),
        (37373,46727,52619,56714,59821,62317,64399,0),
        (37377,46729,52620,56715,59822,62317,64399,0),
        (37379,46731,52621,56715,59822,62318,64400,0),
        (37382,46732,52622,56716,59823,62318,64400,0),
        (37384,46735,52623,56717,59824,62319,64401,0),
        (37388,46736,52624,56718,59824,62319,64401,0),
        (37390,46738,52625,56719,59825,62320,64402,0),
        (37393,46739,52627,56720,59826,62320,64402,0),
        (37397,46742,52628,56721,59826,62321,64403,0),
        (37399,46743,52629,56721,59827,62322,64403,0),
        (37402,46745,52630,56722,59828,62322,64404,0),
        (37404,46747,52631,56723,59828,62323,64404,0),
        (37408,46749,52632,56724,59829,62323,64405,0),
        (37410,46750,52633,56725,59830,62324,64405,0),
        (37413,46752,52635,56726,59831,62324,64405,0),
        (37416,46754,52636,56727,59831,62325,64406,0),
        (37419,46756,52637,56727,59832,62326,64406,0),
        (37421,46757,52638,56728,59833,62326,64407,0),
        (37424,46760,52640,56729,59833,62326,64407,0),
        (37427,46761,52641,56730,59834,62327,64408,0),
        (37430,46763,52642,56731,59835,62328,64408,0),
        (37432,46764,52643,56732,59835,62328,64409,0),
        (37436,46767,52644,56733,59836,62329,64409,0),
        (37439,46768,52645,56733,59836,62329,64410,0),
        (37441,46770,52646,56734,59837,62330,64410,0),
        (37444,46772,52648,56735,59838,62330,64411,0),
        (37447,46774,52649,56736,59838,62331,64411,0),
        (37450,46775,52650,56737,59839,62332,64412,0),
        (37452,46777,52651,56738,59840,62332,64412,0),
        (37456,46779,52652,56739,59841,62333,64412,0),
        (37458,46781,52653,56739,59841,62333,64413,0),
        (37461,46782,52654,56740,59842,62334,64413,0),
        (37463,46784,52656,56741,59843,62334,64414,0),
        (37467,46786,52657,56742,59843,62335,64414,0),
        (37469,46787,52658,56743,59844,62335,64415,0),
        (37472,46789,52659,56744,59845,62336,64415,0),
        (37476,46791,52660,56745,59845,62336,64416,0),
        (37478,46793,52662,56745,59846,62337,64416,0),
        (37481,46794,52663,56746,59847,62338,64417,0),
        (37483,46797,52664,56747,59847,62338,64417,0),
        (37487,46798,52665,56748,59848,62339,64418,0),
        (37489,46800,52666,56749,59849,62339,64418,0),
        (37492,46801,52668,56750,59849,62340,64419,0),
        (37495,46804,52669,56751,59850,62340,64419,0),
        (37498,46805,52670,56751,59851,62341,64420,0),
        (37500,46807,52671,56752,59851,62341,64420,0),
        (37503,46809,52672,56753,59852,62342,64420,0),
        (37506,46811,52673,56754,59853,62342,64421,0),
        (37509,46812,52674,56755,59853,62343,64421,0),
        (37511,46814,52676,56756,59854,62344,64422,0),
        (37515,46816,52677,56757,59855,62344,64422,0),
        (37518,46818,52678,56757,59855,62345,64423,0),
        (37520,46819,52679,56758,59856,62345,64423,0),
        (37522,46821,52680,56759,59857,62346,64424,0),
        (37526,46823,52681,56760,59857,62346,64424,0),
        (37529,46825,52682,56761,59858,62347,64425,0),
        (37531,46826,52684,56762,59859,62347,64425,0),
        (37535,46828,52685,56763,59859,62348,64425,0),
        (37537,46830,52686,56763,59860,62349,64426,0),
        (37540,46832,52687,56764,59861,62349,64427,0),
        (37542,46834,52689,56765,59861,62350,64427,0),
        (37546,46835,52690,56766,59862,62350,64428,0),
        (37548,46837,52691,56767,59863,62351,64428,0),
        (37551,46838,52692,56768,59863,62351,64428,0),
        (37554,46841,52693,56769,59864,62352,64429,0),
        (37557,46842,52694,56769,59865,62353,64429,0),
        (37559,46844,52695,56770,59866,62353,64430,0),
        (37562,46846,52697,56771,59866,62354,64430,0),
        (37566,46848,52698,56772,59867,62354,64431,0),
        (37568,46849,52699,56773,59868,62355,64431,0),
        (37570,46851,52700,56774,59868,62355,64432,0),
        (37574,46853,52701,56775,59869,62356,64432,0),
        (37577,46855,52702,56775,59869,62356,64433,0),
        (37579,46856,52703,56776,59870,62357,64433,0),
        (37582,46858,52705,56777,59871,62357,64433,0),
        (37585,46860,52706,56778,59871,62358,64434,0),
        (37588,46862,52707,56779,59872,62359,64434,0),
        (37590,46863,52708,56780,59873,62359,64435,0),
        (37594,46865,52709,56780,59873,62360,64435,0),
        (37596,46867,52710,56781,59874,62360,64436,0),
        (37599,46869,52712,56782,59875,62361,64436,0),
        (37602,46871,52713,56783,59875,62361,64437,0),
        (37605,46872,52714,56784,59876,62362,64437,0),
        (37607,46874,52715,56785,59877,62362,64438,0),
        (37610,46876,52717,56786,59878,62363,64438,0),
        (37614,46878,52718,56786,59878,62363,64439,0),
        (37616,46879,52719,56787,59879,62364,64439,0),
        (37618,46881,52720,56788,59880,62365,64440,0),
        (37622,46883,52721,56789,59880,62365,64440,0),
        (37625,46885,52722,56790,59881,62366,64441,0),
        (37627,46886,52723,56791,59882,62366,64441,0),
        (37629,46888,52725,56792,59882,62367,64441,0),
        (37633,46890,52726,56792,59883,62367,64442,0),
        (37636,46892,52727,56793,59884,62368,64442,0),
        (37638,46893,52728,56794,59884,62368,64443,0),
        (37642,46895,52729,56795,59885,62369,64443,0),
        (37644,46897,52730,56796,59885,62370,64444,0),
        (37647,46898,52731,56797,59886,62370,64444,0),
        (37649,46901,52733,56798,59887,62371,64445,0),
        (37653,46902,52734,56798,59888,62371,64445,0),
        (37655,46904,52735,56799,59888,62372,64446,0),
        (37658,46905,52736,56800,59889,62372,64446,0),
        (37661,46908,52737,56801,59890,62373,64447,0),
        (37664,46909,52738,56802,59890,62374,64447,0),
        (37666,46911,52739,56803,59891,62374,64448,0),
        (37669,46913,52741,56804,59892,62374,64448,0),
        (37672,46915,52742,56804,59892,62375,64449,0),
        (37675,46916,52743,56805,59893,62376,64449,0),
        (37677,46918,52745,56806,59894,62376,64449,0),
        (37681,46920,52746,56807,59894,62377,64450,0),
        (37683,46922,52747,56808,59895,62377,64450,0),
        (37686,46923,52748,56809,59896,62378,64451,0),
        (37688,46925,52749,56810,59896,62378,64451,0),
        (37692,46927,52750,56810,59897,62379,64452,0),
        (37694,46928,52751,56811,59898,62380,64452,0),
        (37697,46930,52753,56812,59898,62380,64453,0),
        (37701,46932,52754,56813,59899,62381,64453,0),
        (37703,46934,52755,56814,59900,62381,64454,0),
        (37706,46935,52756,56815,59900,62382,64454,0),
        (37708,46938,52757,56816,59901,62382,64455,0),
        (37712,46939,52758,56816,59902,62383,64455,0),
        (37714,46941,52759,56817,59902,62383,64456,0),
        (37717,46942,52761,56818,59903,62384,64456,0),
        (37720,46944,52762,56819,59904,62384,64456,0),
        (37723,46946,52763,56820,59904,62385,64457,0),
        (37725,46948,52764,56821,59905,62386,64457,0),
        (37728,46950,52765,56822,59906,62386,64458,0),
        (37731,46951,52766,56822,59906,62387,64458,0),
        (37734,46953,52767,56823,59907,62387,64459,0),
        (37736,46954,52769,56824,59908,62388,64459,0),
        (37740,46957,52770,56825,59908,62388,64460,0),
        (37742,46958,52771,56826,59909,62389,64460,0),
        (37745,46960,52772,56827,59910,62389,64461,0),
        (37747,46962,52773,56827,59910,62390,64461,0),
        (37751,46964,52774,56828,59911,62390,64462,0),
        (37753,46965,52776,56829,59912,62391,64462,0),
        (37756,46967,52777,56830,59912,62392,64462,0),
        (37759,46969,52778,56831,59913,62392,64463,0),
        (37762,46970,52779,56832,59914,62393,64463,0),
        (37764,46972,52780,56833,59914,62393,64464,0),
        (37767,46974,52782,56833,59915,62394,64464,0),
        (37770,46976,52783,56834,59916,62394,64465,0),
        (37773,46977,52784,56835,59916,62395,64465,0),
        (37775,46979,52785,56836,59917,62395,64466,0),
        (37779,46981,52786,56837,59918,62396,64466,0),
        (37781,46983,52787,56838,59918,62397,64467,0),
        (37784,46984,52788,56839,59919,62397,64467,0),
        (37786,46987,52790,56839,59920,62398,64468,0),
        (37790,46988,52791,56840,59920,62398,64468,0),
        (37792,46990,52792,56841,59921,62399,64469,0),
        (37795,46991,52793,56842,59922,62399,64469,0),
        (37799,46993,52794,56843,59922,62400,64469,0),
        (37801,46995,52795,56843,59923,62400,64470,0),
        (37803,46996,52796,56845,59924,62401,64470,0),
        (37806,46999,52798,56845,59924,62401,64471,0),
        (37809,47000,52799,56846,59925,62402,64471,0),
        (37812,47002,52800,56847,59926,62403,64472,0),
        (37814,47003,52801,56848,59926,62403,64472,0),
        (37818,47006,52802,56849,59927,62404,64473,0),
        (37820,47007,52803,56849,59928,62404,64473,0),
        (37823,47009,52804,56851,59928,62405,64474,0),
        (37825,47011,52806,56851,59929,62405,64474,0),
        (37829,47012,52807,56852,59930,62406,64475,0),
        (37831,47014,52808,56853,59931,62406,64475,0),
        (37834,47016,52809,56854,59931,62407,64476,0),
        (37838,47018,52810,56855,59932,62407,64476,0),
        (37840,47019,52811,56855,59932,62408,64477,0),
        (37842,47021,52812,56856,59933,62409,64477,0),
        (37845,47023,52814,56857,59934,62409,64477,0),
        (37849,47025,52815,56858,59934,62410,64478,0),
        (37851,47026,52816,56859,59935,62410,64478,0),
        (37853,47028,52818,56860,59936,62411,64479,0),
        (37857,47030,52819,56861,59936,62411,64479,0),
        (37860,47032,52820,56861,59937,62412,64480,0),
        (37862,47033,52821,56862,59938,62412,64480,0),
        (37864,47035,52822,56863,59938,62413,64481,0),
        (37868,47037,52823,56864,59939,62413,64481,0),
        (37870,47038,52824,56865,59940,62414,64482,0),
        (37873,47040,52826,56866,59940,62415,64482,0),
        (37877,47042,52827,56866,59941,62415,64482,0),
        (37879,47044,52828,56867,59942,62416,64483,0),
        (37881,47045,52829,56868,59942,62416,64483,0),
        (37884,47047,52830,56869,59943,62417,64484,0),
        (37888,47049,52831,56870,59944,62417,64484,0),
        (37890,47051,52832,56871,59945,62418,64485,0),
        (37892,47052,52834,56872,59945,62418,64485,0),
        (37896,47054,52835,56872,59946,62419,64486,0),
        (37899,47056,52836,56873,59946,62420,64486,0),
        (37901,47057,52837,56874,59947,62420,64487,0),
        (37903,47060,52838,56875,59948,62421,64487,0),
        (37907,47061,52839,56876,59948,62421,64488,0),
        (37909,47063,52840,56877,59949,62422,64488,0),
        (37912,47064,52842,56878,59950,62422,64489,0),
        (37916,47066,52843,56878,59950,62423,64489,0),
        (37918,47068,52844,56879,59951,62424,64490,0),
        (37920,47070,52845,56880,59952,62424,64490,0),
        (37923,47072,52846,56881,59952,62424,64490,0),
        (37927,47073,52847,56882,59953,62425,64491,0),
        (37929,47075,52848,56882,59954,62426,64491,0),
        (37931,47076,52850,56884,59954,62426,64492,0),
        (37935,47079,52851,56884,59955,62427,64492,0),
        (37937,47080,52852,56885,59956,62427,64493,0),
        (37940,47082,52853,56886,59956,62428,64493,0),
        (37942,47084,52854,56887,59957,62428,64494,0),
        (37946,47085,52855,56888,59958,62429,64494,0),
        (37948,47087,52856,56888,59959,62430,64495,0),
        (37951,47089,52858,56889,59959,62430,64495,0),
        (37954,47091,52859,56890,59960,62430,64495,0),
        (37957,47092,52860,56891,59960,62431,64496,0),
        (37959,47094,52861,56892,59961,62432,64496,0),
        (37962,47096,52862,56893,59962,62432,64497,0),
        (37965,47098,52863,56894,59962,62433,64497,0),
        (37968,47099,52864,56894,59963,62433,64498,0),
        (37970,47101,52866,56895,59964,62434,64498,0),
        (37974,47103,52867,56896,59964,62434,64499,0),
        (37976,47104,52868,56897,59965,62435,64499,0),
        (37979,47106,52869,56898,59966,62436,64500,0),
        (37981,47108,52870,56899,59966,62436,64500,0),
        (37985,47110,52871,56899,59967,62436,64501,0),
        (37987,47111,52872,56900,59968,62437,64501,0),
        (37990,47113,52874,56901,59968,62438,64502,0),
        (37993,47115,52875,56902,59969,62438,64502,0),
        (37996,47117,52876,56903,59970,62439,64503,0),
        (37998,47118,52877,56904,59970,62439,64503,0),
        (38001,47120,52878,56905,59971,62440,64503,0),
        (38004,47122,52879,56905,59972,62440,64504,0),
        (38007,47123,52880,56906,59973,62441,64504,0),
        (38009,47125,52882,56907,59973,62441,64505,0),
        (38013,47127,52883,56908,59974,62442,64505,0),
        (38015,47129,52884,56909,59974,62443,64506,0),
        (38018,47130,52885,56910,59975,62443,64506,0),
        (38020,47132,52887,56911,59976,62444,64507,0),
        (38024,47134,52888,56911,59976,62444,64507,0),
        (38026,47135,52889,56912,59977,62445,64508,0),
        (38029,47137,52890,56913,59978,62445,64508,0),
        (38032,47139,52891,56914,59978,62446,64508,0),
        (38035,47141,52892,56915,59979,62447,64509,0),
        (38037,47142,52893,56916,59980,62447,64509,0),
        (38039,47145,52895,56916,59980,62447,64510,0),
        (38043,47146,52896,56917,59981,62448,64510,0),
        (38046,47148,52897,56918,59982,62449,64511,0),
        (38048,47149,52898,56919,59982,62449,64511,0),
        (38052,47151,52899,56920,59983,62450,64512,0),
        (38054,47153,52900,56921,59984,62450,64512,0),
        (38056,47154,52901,56922,59984,62451,64513,0),
        (38059,47157,52903,56922,59985,62451,64513,0),
        (38062,47158,52904,56923,59986,62452,64514,0),
        (38065,47160,52905,56924,59986,62453,64514,0),
        (38067,47161,52906,56925,59987,62453,64515,0),
        (38071,47163,52907,56926,59988,62453,64515,0),
        (38073,47165,52908,56926,59988,62454,64516,0),
        (38076,47166,52909,56928,59989,62455,64516,0),
        (38078,47169,52911,56928,59990,62455,64516,0),
        (38082,47170,52912,56929,59990,62456,64517,0),
        (38084,47172,52913,56930,59991,62456,64517,0),
        (38087,47173,52914,56931,59992,62457,64518,0),
        (38090,47175,52915,56932,59992,62457,64518,0),
        (38093,47177,52916,56932,59993,62458,64519,0),
        (38095,47178,52917,56933,59994,62458,64519,0),
        (38098,47181,52919,56934,59994,62459,64520,0),
        (38101,47182,52920,56935,59995,62459,64520,0),
        (38104,47184,52921,56936,59996,62460,64521,0),
        (38106,47185,52922,56937,59996,62461,64521,0),
        (38110,47188,52923,56938,59997,62461,64521,0),
        (38112,47189,52924,56938,59998,62462,64522,0),
        (38115,47191,52925,56939,59998,62462,64522,0),
        (38117,47193,52927,56940,59999,62463,64523,0),
        (38121,47194,52928,56941,60000,62463,64523,0),
        (38123,47196,52929,56942,60000,62464,64524,0),
        (38125,47197,52930,56943,60001,62464,64524,0),
        (38129,47200,52931,56943,60002,62465,64525,0),
        (38131,47201,52932,56944,60002,62466,64525,0),
        (38134,47203,52933,56945,60003,62466,64526,0),
        (38136,47205,52935,56946,60004,62467,64526,0),
        (38140,47206,52936,56947,60004,62467,64527,0),
        (38142,47208,52937,56948,60005,62468,64527,0),
        (38145,47209,52938,56949,60006,62468,64528,0),
        (38148,47212,52939,56949,60006,62469,64528,0),
        (38151,47213,52940,56950,60007,62469,64529,0),
        (38153,47215,52941,56951,60008,62470,64529,0),
        (38156,47217,52943,56952,60008,62470,64529,0),
        (38159,47218,52944,56953,60009,62471,64530,0),
        (38162,47220,52945,56953,60010,62472,64530,0),
        (38164,47221,52946,56955,60010,62472,64531,0),
        (38168,47224,52947,56955,60011,62473,64531,0),
        (38170,47225,52948,56956,60011,62473,64532,0),
        (38173,47227,52949,56957,60012,62474,64532,0),
        (38175,47229,52951,56958,60013,62474,64533,0),
        (38179,47230,52952,56959,60013,62475,64533,0),
        (38181,47232,52953,56959,60014,62475,64534,0),
        (38183,47233,52954,56960,60015,62476,64534,0),
        (38187,47236,52955,56961,60016,62476,64534,0),
        (38189,47237,52956,56962,60016,62477,64535,0),
        (38192,47239,52957,56963,60017,62478,64535,0),
        (38194,47241,52959,56964,60018,62478,64536,0),
        (38198,47242,52960,56964,60018,62479,64536,0),
        (38200,47244,52961,56965,60019,62479,64537,0),
        (38203,47245,52962,56966,60020,62480,64537,0),
        (38206,47248,52963,56967,60020,62480,64538,0),
        (38209,47249,52964,56968,60021,62481,64538,0),
        (38211,47251,52965,56969,60022,62481,64539,0),
        (38214,47253,52967,56970,60022,62482,64539,0),
        (38217,47254,52968,56970,60023,62482,64540,0),
        (38220,47256,52969,56971,60024,62483,64540,0),
        (38222,47257,52970,56972,60024,62484,64541,0),
        (38226,47260,52971,56973,60025,62484,64541,0),
        (38228,47261,52972,56974,60025,62485,64542,0),
        (38230,47263,52973,56975,60026,62485,64542,0),
        (38233,47265,52975,56976,60027,62486,64542,0),
        (38236,47266,52976,56976,60027,62486,64543,0),
        (38239,47268,52977,56977,60028,62487,64543,0),
        (38241,47269,52978,56978,60029,62487,64544,0),
        (38245,47272,52979,56979,60029,62488,64544,0),
        (38247,47273,52980,56980,60030,62489,64545,0),
        (38250,47275,52981,56981,60031,62489,64545,0),
        (38252,47277,52983,56981,60031,62490,64546,0),
        (38256,47278,52984,56982,60032,62490,64546,0),
        (38258,47280,52985,56983,60033,62491,64547,0),
        (38261,47281,52986,56984,60033,62491,64547,0),
        (38264,47284,52987,56985,60034,62492,64547,0),
        (38267,47285,52988,56985,60035,62492,64548,0),
        (38269,47287,52989,56987,60036,62493,64548,0),
        (38271,47289,52991,56987,60036,62493,64549,0),
        (38275,47290,52992,56988,60037,62494,64549,0),
        (38277,47292,52993,56989,60038,62495,64550,0),
        (38280,47293,52994,56990,60038,62495,64550,0),
        (38283,47296,52995,56991,60039,62496,64551,0),
        (38286,47297,52996,56991,60039,62496,64551,0),
        (38288,47299,52997,56992,60040,62497,64552,0),
        (38291,47301,52999,56993,60041,62497,64552,0),
        (38294,47302,53000,56994,60041,62498,64553,0),
        (38297,47304,53001,56995,60042,62498,64553,0),
        (38299,47305,53002,56996,60043,62499,64553,0),
        (38303,47308,53003,56996,60043,62499,64554,0),
        (38305,47309,53004,56997,60044,62500,64554,0),
        (38307,47311,53005,56998,60045,62501,64555,0),
        (38310,47313,53007,56999,60045,62501,64555,0),
        (38313,47314,53008,57000,60046,62501,64556,0),
        (38316,47316,53009,57001,60047,62502,64556,0),
        (38318,47317,53010,57002,60047,62503,64557,0),
        (38322,47320,53011,57002,60048,62503,64557,0),
        (38324,47321,53012,57003,60049,62504,64558,0),
        (38327,47323,53013,57004,60049,62504,64558,0),
        (38329,47325,53015,57005,60050,62505,64559,0),
        (38333,47326,53016,57006,60051,62505,64559,0),
        (38335,47328,53017,57006,60051,62506,64560,0),
        (38337,47329,53018,57007,60052,62506,64560,0),
        (38341,47331,53019,57008,60053,62507,64560,0),
        (38343,47333,53020,57009,60053,62508,64561,0),
        (38346,47334,53021,57010,60054,62508,64561,0),
        (38348,47337,53023,57011,60055,62509,64562,0),
        (38352,47338,53024,57012,60055,62509,64562,0),
        (38354,47340,53025,57012,60056,62510,64563,0),
        (38357,47341,53026,57013,60057,62510,64563,0),
        (38360,47343,53027,57014,60057,62511,64564,0),
        (38363,47345,53028,57015,60058,62511,64564,0),
        (38365,47346,53029,57016,60059,62512,64565,0),
        (38369,47349,53030,57017,60059,62512,64565,0),
        (38371,47350,53031,57017,60060,62513,64566,0),
        (38373,47352,53032,57018,60061,62514,64566,0),
        (38376,47354,53034,57019,60061,62514,64566,0),
        (38379,47355,53035,57020,60062,62515,64567,0),
        (38382,47357,53036,57021,60063,62515,64567,0),
        (38384,47358,53037,57022,60063,62516,64568,0),
        (38388,47361,53038,57023,60064,62516,64568,0),
        (38390,47362,53039,57023,60064,62517,64569,0),
        (38393,47364,53040,57024,60065,62517,64569,0),
        (38395,47366,53042,57025,60066,62518,64570,0),
        (38399,47367,53043,57026,60066,62518,64570,0),
        (38401,47369,53044,57027,60067,62519,64571,0),
        (38403,47370,53045,57028,60068,62520,64571,0),
        (38407,47372,53046,57028,60069,62520,64571,0),
        (38409,47374,53047,57029,60069,62521,64572,0),
        (38412,47375,53048,57030,60070,62521,64573,0),
        (38414,47378,53050,57031,60071,62522,64573,0),
        (38418,47379,53051,57032,60071,62522,64574,0),
        (38420,47381,53052,57032,60072,62523,64574,0),
        (38423,47382,53053,57034,60073,62523,64574,0),
        (38426,47384,53054,57034,60073,62524,64575,0),
        (38429,47386,53055,57035,60074,62525,64575,0),
        (38431,47387,53056,57036,60075,62525,64576,0),
        (38433,47390,53058,57037,60075,62526,64576,0),
        (38437,47391,53059,57038,60076,62526,64577,0),
        (38439,47393,53060,57038,60077,62527,64577,0),
        (38442,47394,53061,57039,60077,62527,64578,0),
        (38445,47396,53062,57040,60078,62528,64578,0),
        (38448,47398,53063,57041,60078,62528,64579,0),
        (38450,47399,53064,57042,60079,62529,64579,0),
        (38452,47401,53066,57043,60080,62529,64579,0),
        (38456,47403,53067,57043,60080,62530,64580,0),
        (38458,47404,53068,57044,60081,62531,64580,0),
        (38461,47406,53069,57045,60082,62531,64581,0),
        (38464,47408,53070,57046,60082,62531,64581,0),
        (38467,47410,53071,57047,60083,62532,64582,0),
        (38469,47411,53072,57048,60084,62533,64582,0),
        (38472,47413,53074,57049,60084,62533,64583,0),
        (38475,47415,53075,57049,60085,62534,64583,0),
        (38478,47416,53076,57050,60086,62534,64584,0),
        (38480,47418,53077,57051,60086,62535,64584,0),
        (38484,47420,53078,57052,60087,62535,64584,0),
        (38486,47422,53079,57053,60088,62536,64585,0),
        (38488,47423,53080,57054,60088,62536,64585,0),
        (38491,47425,53082,57054,60089,62537,64586,0),
        (38494,47427,53083,57055,60090,62537,64586,0),
        (38497,47428,53084,57056,60090,62538,64587,0),
        (38499,47430,53085,57057,60091,62539,64587,0),
        (38503,47432,53086,57058,60092,62539,64588,0),
        (38505,47433,53087,57058,60092,62540,64588,0),
        (38507,47435,53088,57059,60093,62540,64589,0),
        (38510,47437,53090,57060,60094,62541,64589,0),
        (38513,47439,53091,57061,60094,62541,64590,0),
        (38516,47440,53092,57062,60095,62542,64590,0),
        (38518,47442,53093,57063,60096,62542,64590,0),
        (38522,47444,53094,57064,60096,62543,64591,0),
        (38524,47445,53095,57064,60097,62544,64591,0),
        (38526,47447,53096,57065,60098,62544,64592,0),
        (38529,47449,53097,57066,60098,62545,64592,0),
        (38532,47450,53098,57067,60099,62545,64593,0),
        (38535,47452,53099,57068,60100,62546,64593,0),
        (38537,47453,53101,57069,60100,62546,64594,0),
        (38541,47456,53102,57069,60101,62547,64594,0),
        (38543,47457,53103,57070,60101,62547,64595,0),
        (38546,47459,53104,57071,60102,62548,64595,0),
        (38548,47461,53105,57072,60103,62548,64596,0),
        (38552,47462,53106,57073,60103,62549,64596,0),
        (38554,47464,53107,57073,60104,62550,64597,0),
        (38556,47465,53109,57074,60105,62550,64597,0),
        (38560,47467,53110,57075,60105,62550,64597,0),
        (38562,47469,53111,57076,60106,62551,64598,0),
        (38565,47470,53112,57077,60107,62552,64598,0),
        (38567,47473,53113,57078,60107,62552,64599,0),
        (38571,47474,53114,57078,60108,62553,64599,0),
        (38573,47476,53115,57079,60109,62553,64600,0),
        (38575,47477,53117,57080,60109,62554,64600,0),
        (38579,47479,53118,57081,60110,62554,64601,0),
        (38581,47481,53119,57082,60111,62555,64601,0),
        (38584,47482,53120,57083,60111,62555,64602,0),
        (38586,47484,53121,57084,60112,62556,64602,0),
        (38590,47486,53122,57084,60113,62556,64603,0),
        (38592,47487,53123,57085,60113,62557,64603,0),
        (38594,47489,53125,57086,60114,62558,64603,0),
        (38598,47491,53126,57087,60115,62558,64604,0),
        (38600,47493,53127,57088,60115,62559,64604,0),
        (38603,47494,53128,57089,60116,62559,64605,0),
        (38605,47496,53129,57089,60117,62560,64605,0),
        (38609,47498,53130,57090,60117,62560,64606,0),
        (38611,47499,53131,57091,60118,62561,64606,0),
        (38613,47501,53133,57092,60119,62561,64607,0),
        (38617,47503,53134,57093,60119,62562,64607,0),
        (38619,47504,53134,57093,60120,62563,64608,0),
        (38622,47506,53135,57095,60121,62563,64608,0),
        (38624,47508,53137,57095,60121,62564,64608,0),
        (38628,47510,53138,57096,60122,62564,64609,0),
        (38630,47511,53139,57097,60123,62565,64609,0),
        (38632,47512,53140,57098,60123,62565,64610,0),
        (38636,47515,53141,57099,60124,62566,64610,0),
        (38638,47516,53142,57099,60124,62566,64611,0),
        (38641,47518,53143,57100,60125,62567,64611,0),
        (38643,47520,53145,57101,60126,62567,64612,0),
        (38647,47521,53146,57102,60126,62568,64612,0),
        (38649,47523,53147,57103,60127,62569,64613,0),
        (38651,47524,53148,57104,60128,62569,64613,0),
        (38655,47526,53149,57104,60128,62569,64613,0),
        (38657,47528,53150,57105,60129,62570,64614,0),
        (38660,47529,53151,57106,60130,62571,64614,0),
        (38662,47532,53153,57107,60130,62571,64615,0),
        (38666,47533,53154,57108,60131,62572,64615,0),
        (38668,47535,53155,57108,60132,62572,64616,0),
        (38670,47536,53156,57109,60132,62573,64616,0),
        (38674,47538,53157,57110,60133,62573,64617,0),
        (38676,47540,53158,57111,60134,62574,64617,0),
        (38679,47541,53159,57112,60134,62574,64618,0),
        (38681,47543,53161,57113,60135,62575,64618,0),
        (38685,47545,53162,57113,60136,62575,64619,0),
        (38687,47546,53163,57114,60137,62576,64619,0),
        (38689,47548,53164,57115,60137,62577,64620,0),
        (38693,47550,53165,57116,60138,62577,64620,0),
        (38695,47552,53166,57117,60138,62578,64621,0),
        (38698,47553,53167,57118,60139,62578,64621,0),
        (38700,47555,53168,57119,60140,62579,64621,0),
        (38704,47557,53169,57119,60140,62579,64622,0),
        (38706,47558,53170,57120,60141,62580,64622,0),
        (38708,47560,53172,57121,60142,62580,64623,0),
        (38712,47562,53173,57122,60142,62581,64623,0),
        (38714,47563,53174,57123,60143,62582,64624,0),
        (38717,47565,53175,57124,60144,62582,64624,0),
        (38719,47567,53176,57124,60144,62582,64625,0),
        (38723,47568,53177,57125,60145,62583,64625,0),
        (38725,47570,53178,57126,60146,62584,64626,0),
        (38727,47571,53180,57127,60146,62584,64626,0),
        (38731,47574,53181,57128,60147,62585,64626,0),
        (38733,47575,53182,57128,60147,62585,64627,0),
        (38736,47576,53183,57130,60148,62586,64627,0),
        (38738,47579,53184,57130,60149,62586,64628,0),
        (38742,47580,53185,57131,60149,62587,64628,0),
        (38744,47582,53186,57132,60150,62587,64629,0),
        (38746,47583,53188,57133,60151,62588,64629,0),
        (38750,47585,53189,57133,60151,62588,64630,0),
        (38752,47587,53190,57134,60152,62589,64630,0),
        (38755,47588,53191,57135,60153,62590,64631,0),
        (38757,47590,53192,57136,60153,62590,64631,0),
        (38760,47592,53193,57137,60154,62591,64632,0),
        (38763,47593,53194,57137,60155,62591,64632,0),
        (38765,47595,53196,57139,60155,62592,64632,0),
        (38769,47597,53197,57139,60156,62592,64633,0),
        (38771,47598,53197,57140,60157,62593,64633,0),
        (38773,47600,53198,57141,60157,62593,64634,0),
        (38776,47602,53200,57142,60158,62594,64634,0),
        (38779,47604,53201,57143,60159,62594,64635,0),
        (38782,47605,53202,57143,60159,62595,64635,0),
        (38784,47607,53203,57144,60160,62596,64636,0),
        (38788,47609,53204,57145,60161,62596,64636,0),
        (38790,47610,53205,57146,60161,62597,64637,0),
        (38792,47612,53206,57147,60162,62597,64637,0),
        (38795,47614,53208,57148,60163,62598,64637,0),
        (38798,47615,53209,57148,60163,62598,64638,0),
        (38801,47617,53210,57149,60164,62599,64638,0),
        (38803,47618,53211,57150,60165,62599,64639,0),
        (38807,47620,53212,57151,60165,62600,64639,0),
        (38809,47622,53213,57152,60166,62600,64640,0),
        (38811,47623,53214,57153,60167,62601,64640,0),
        (38814,47626,53216,57153,60167,62601,64641,0),
        (38817,47627,53217,57154,60168,62602,64641,0),
        (38820,47629,53218,57155,60169,62603,64642,0),
        (38822,47630,53219,57156,60169,62603,64642,0),
        (38825,47632,53220,57157,60170,62604,64642,0),
        (38828,47634,53221,57157,60170,62604,64643,0),
        (38830,47635,53222,57159,60171,62605,64643,0),
        (38833,47637,53223,57159,60172,62605,64644,0),
        (38836,47639,53224,57160,60172,62606,64644,0),
        (38838,47640,53225,57161,60173,62606,64645,0),
        (38841,47642,53227,57162,60174,62607,64645,0),
        (38844,47644,53228,57163,60174,62607,64646,0),
        (38847,47645,53229,57163,60175,62608,64646,0),
        (38849,47647,53230,57164,60176,62609,64647,0),
        (38851,47649,53231,57165,60176,62609,64647,0),
        (38855,47650,53232,57166,60177,62609,64648,0),
        (38857,47652,53233,57167,60178,62610,64648,0),
        (38860,47653,53235,57168,60178,62611,64648,0),
        (38863,47656,53236,57168,60179,62611,64649,0),
        (38866,47657,53237,57169,60180,62612,64649,0),
        (38868,47658,53238,57170,60180,62612,64650,0),
        (38870,47661,53239,57171,60181,62613,64650,0),
        (38874,47662,53240,57172,60182,62613,64651,0),
        (38876,47664,53241,57172,60182,62614,64651,0),
        (38878,47665,53243,57173,60183,62614,64652,0),
        (38882,47667,53244,57174,60184,62615,64652,0),
        (38884,47669,53245,57175,60184,62616,64653,0),
        (38887,47670,53246,57176,60185,62616,64653,0),
        (38889,47672,53247,57177,60186,62617,64654,0),
        (38893,47674,53248,57177,60186,62617,64654,0),
        (38895,47675,53249,57178,60187,62618,64655,0),
        (38897,47677,53250,57179,60188,62618,64655,0),
        (38901,47679,53251,57180,60188,62619,64655,0),
        (38903,47680,53252,57181,60189,62619,64656,0),
        (38906,47682,53253,57182,60190,62620,64656,0),
        (38908,47684,53255,57182,60190,62620,64657,0),
        (38911,47685,53256,57183,60191,62621,64657,0),
        (38914,47687,53257,57184,60192,62621,64658,0),
        (38916,47688,53258,57185,60192,62622,64658,0),
        (38920,47691,53259,57186,60193,62622,64659,0),
        (38922,47692,53260,57186,60193,62623,64659,0),
        (38924,47693,53261,57188,60194,62624,64660,0),
        (38927,47696,53263,57188,60195,62624,64660,0),
        (38930,47697,53264,57189,60195,62625,64661,0),
        (38933,47699,53265,57190,60196,62625,64661,0),
        (38935,47700,53266,57191,60197,62626,64661,0),
        (38938,47702,53267,57192,60197,62626,64662,0),
        (38941,47704,53268,57192,60198,62627,64662,0),
        (38943,47705,53269,57193,60199,62627,64663,0),
        (38946,47707,53270,57194,60199,62628,64663,0),
        (38949,47709,53271,57195,60200,62628,64664,0),
        (38951,47710,53272,57196,60201,62629,64664,0),
        (38954,47712,53274,57197,60201,62630,64665,0),
        (38957,47714,53275,57197,60202,62630,64665,0),
        (38960,47715,53276,57198,60202,62631,64666,0),
        (38962,47717,53277,57199,60203,62631,64666,0),
        (38964,47719,53278,57200,60204,62632,64666,0),
        (38968,47720,53279,57201,60204,62632,64667,0),
        (38970,47722,53280,57201,60205,62633,64667,0),
        (38973,47723,53282,57202,60206,62633,64668,0),
        (38976,47725,53283,57203,60206,62634,64668,0),
        (38978,47727,53284,57204,60207,62634,64669,0),
        (38981,47728,53285,57205,60208,62635,64669,0),
        (38983,47731,53286,57206,60208,62635,64670,0),
        (38987,47732,53287,57206,60209,62636,64670,0),
        (38989,47733,53288,57207,60210,62637,64671,0),
        (38991,47735,53289,57208,60210,62637,64671,0),
        (38995,47737,53290,57209,60211,62638,64671,0),
        (38997,47739,53291,57210,60212,62638,64672,0),
        (38999,47740,53292,57211,60212,62639,64672,0),
        (39002,47742,53294,57211,60213,62639,64673,0),
        (39005,47744,53295,57212,60214,62640,64673,0),
        (39008,47745,53296,57213,60214,62640,64674,0),
        (39010,47747,53297,57214,60215,62641,64674,0),
        (39014,47749,53298,57215,60216,62641,64675,0),
        (39016,47750,53299,57215,60216,62642,64675,0),
        (39018,47752,53300,57216,60217,62642,64676,0),
        (39021,47754,53302,57217,60218,62643,64676,0),
        (39024,47755,53303,57218,60218,62643,64677,0),
        (39026,47757,53304,57219,60219,62644,64677,0),
        (39029,47758,53305,57220,60220,62645,64677,0),
        (39032,47760,53306,57220,60220,62645,64678,0),
        (39035,47762,53307,57221,60221,62646,64678,0),
        (39037,47763,53308,57222,60222,62646,64679,0),
        (39039,47765,53309,57223,60222,62647,64679,0),
        (39043,47767,53310,57224,60223,62647,64680,0),
        (39045,47768,53311,57224,60224,62648,64680,0),
        (39048,47770,53313,57225,60224,62648,64681,0),
        (39051,47772,53314,57226,60225,62649,64681,0),
        (39053,47773,53315,57227,60225,62650,64682,0),
        (39056,47775,53316,57228,60226,62650,64682,0),
        (39058,47777,53317,57229,60227,62651,64682,0),
        (39062,47778,53318,57229,60227,62651,64683,0),
        (39064,47780,53319,57230,60228,62652,64683,0),
        (39066,47781,53321,57231,60229,62652,64684,0),
        (39070,47784,53322,57232,60229,62653,64684,0),
        (39072,47785,53323,57233,60230,62653,64685,0),
        (39074,47786,53324,57234,60231,62654,64685,0),
        (39077,47789,53325,57235,60231,62654,64686,0),
        (39080,47790,53326,57235,60232,62655,64686,0),
        (39083,47791,53327,57236,60233,62655,64687,0),
        (39085,47793,53328,57237,60233,62656,64687,0),
        (39088,47795,53329,57238,60234,62656,64687,0),
        (39091,47797,53330,57238,60234,62657,64688,0),
        (39093,47798,53331,57240,60235,62658,64688,0),
        (39095,47800,53333,57240,60236,62658,64689,0),
        (39099,47802,53334,57241,60236,62659,64689,0),
        (39101,47803,53335,57242,60237,62659,64690,0),
        (39104,47805,53336,57243,60238,62660,64690,0),
        (39107,47807,53337,57244,60238,62660,64691,0),
        (39109,47808,53338,57244,60239,62661,64691,0),
        (39112,47810,53340,57245,60240,62661,64692,0),
        (39115,47812,53341,57246,60240,62662,64692,0),
        (39118,47813,53342,57247,60241,62663,64693,0),
        (39120,47815,53343,57248,60242,62663,64693,0),
        (39122,47817,53344,57249,60242,62663,64693,0),
        (39126,47818,53345,57249,60243,62664,64694,0),
        (39128,47820,53346,57250,60244,62665,64694,0),
        (39130,47821,53347,57251,60244,62665,64695,0),
        (39134,47823,53348,57252,60245,62666,64695,0),
        (39136,47825,53349,57253,60246,62666,64696,0),
        (39139,47826,53350,57254,60246,62667,64696,0),
        (39141,47828,53352,57254,60247,62667,64697,0),
        (39144,47830,53353,57255,60248,62668,64697,0),
        (39147,47831,53354,57256,60248,62668,64698,0),
        (39149,47833,53355,57257,60249,62669,64698,0),
        (39153,47835,53356,57258,60250,62669,64698,0),
        (39155,47836,53357,57258,60250,62670,64699,0),
        (39157,47838,53358,57259,60251,62671,64699,0),
        (39160,47840,53360,57260,60252,62671,64700,0),
        (39163,47841,53360,57261,60252,62671,64700,0),
        (39165,47843,53361,57262,60253,62672,64701,0),
        (39168,47844,53363,57263,60254,62673,64701,0),
        (39171,47846,53364,57263,60254,62673,64702,0),
        (39174,47848,53365,57264,60255,62674,64702,0),
        (39176,47849,53366,57265,60256,62674,64703,0),
        (39178,47851,53367,57266,60256,62675,64703,0),
        (39182,47853,53368,57267,60257,62675,64704,0),
        (39184,47854,53369,57267,60257,62676,64704,0),
        (39186,47856,53371,57268,60258,62676,64704,0),
        (39190,47858,53372,57269,60259,62677,64705,0),
        (39192,47859,53373,57270,60259,62678,64705,0),
        (39195,47861,53374,57271,60260,62678,64706,0),
        (39197,47863,53375,57272,60261,62679,64706,0),
        (39200,47864,53376,57272,60261,62679,64707,0),
        (39203,47866,53377,57273,60262,62680,64707,0),
        (39205,47867,53378,57274,60263,62680,64708,0),
        (39209,47869,53379,57275,60263,62681,64708,0),
        (39211,47871,53380,57276,60264,62681,64709,0),
        (39213,47872,53381,57277,60265,62682,64709,0),
        (39215,47874,53383,57277,60265,62682,64709,0),
        (39219,47876,53384,57278,60266,62683,64710,0),
        (39221,47877,53385,57279,60267,62683,64710,0),
        (39224,47879,53386,57280,60267,62684,64711,0),
        (39227,47881,53387,57281,60268,62684,64711,0),
        (39229,47882,53388,57281,60268,62685,64712,0),
        (39232,47884,53389,57282,60269,62686,64712,0),
        (39234,47886,53391,57283,60270,62686,64713,0),
        (39238,47887,53391,57284,60270,62686,64713,0),
        (39240,47889,53392,57285,60271,62687,64714,0),
        (39242,47890,53394,57286,60272,62688,64714,0),
        (39246,47892,53395,57286,60272,62688,64714,0),
        (39248,47894,53396,57287,60273,62689,64715,0),
        (39250,47895,53397,57288,60274,62689,64715,0),
        (39253,47897,53398,57289,60274,62690,64716,0),
        (39256,47899,53399,57290,60275,62690,64716,0),
        (39258,47900,53400,57290,60276,62691,64717,0),
        (39261,47902,53402,57291,60276,62691,64717,0),
        (39264,47904,53403,57292,60277,62692,64718,0),
        (39267,47905,53404,57293,60277,62693,64718,0),
        (39269,47907,53405,57294,60278,62693,64719,0),
        (39271,47909,53406,57295,60279,62694,64719,0),
        (39275,47910,53407,57295,60279,62694,64720,0),
        (39277,47912,53408,57296,60280,62695,64720,0),
        (39279,47913,53409,57297,60281,62695,64720,0),
        (39283,47915,53410,57298,60281,62696,64721,0),
        (39285,47917,53411,57299,60282,62696,64721,0),
        (39287,47918,53412,57300,60283,62697,64722,0),
        (39290,47920,53414,57300,60283,62697,64722,0),
        (39293,47922,53415,57301,60284,62698,64723,0),
        (39296,47923,53416,57302,60285,62698,64723,0),
        (39298,47925,53417,57303,60285,62699,64724,0),
        (39301,47927,53418,57304,60286,62699,64724,0),
        (39304,47928,53419,57304,60286,62700,64725,0),
        (39306,47930,53420,57305,60287,62701,64725,0),
        (39308,47932,53421,57306,60288,62701,64725,0),
        (39312,47933,53422,57307,60288,62702,64726,0),
        (39314,47935,53423,57308,60289,62702,64726,0),
        (39316,47936,53425,57309,60290,62703,64727,0),
        (39320,47938,53426,57309,60290,62703,64727,0),
        (39322,47940,53427,57310,60291,62704,64728,0),
        (39325,47941,53428,57311,60292,62704,64728,0),
        (39327,47943,53429,57312,60292,62705,64729,0),
        (39330,47945,53430,57313,60293,62705,64729,0),
        (39333,47946,53431,57313,60294,62706,64730,0),
        (39335,47948,53433,57314,60294,62706,64730,0),
        (39338,47950,53434,57315,60295,62707,64730,0),
        (39341,47951,53434,57316,60296,62708,64731,0),
        (39343,47953,53435,57317,60296,62708,64731,0),
        (39345,47955,53437,57318,60297,62709,64732,0),
        (39349,47956,53438,57318,60298,62709,64732,0),
        (39351,47958,53439,57319,60298,62710,64733,0),
        (39353,47959,53440,57320,60299,62710,64733,0),
        (39357,47961,53441,57321,60300,62711,64734,0),
        (39359,47963,53442,57321,60300,62711,64734,0),
        (39362,47964,53443,57323,60301,62712,64735,0),
        (39364,47966,53445,57323,60302,62712,64735,0),
        (39367,47968,53446,57324,60302,62713,64736,0),
        (39370,47969,53447,57325,60303,62713,64736,0),
        (39372,47971,53448,57326,60304,62714,64736,0),
        (39375,47973,53449,57327,60304,62714,64737,0),
        (39378,47974,53450,57327,60305,62715,64737,0),
        (39380,47976,53451,57328,60306,62716,64738,0),
        (39382,47978,53452,57329,60306,62716,64738,0),
        (39386,47979,53453,57330,60307,62717,64739,0),
        (39388,47981,53454,57330,60307,62717,64739,0),
        (39390,47982,53456,57332,60308,62718,64740,0),
        (39394,47984,53457,57332,60309,62718,64740,0),
        (39396,47986,53458,57333,60309,62719,64741,0),
        (39399,47987,53459,57334,60310,62719,64741,0),
        (39401,47989,53460,57335,60311,62720,64741,0),
        (39404,47991,53461,57335,60311,62720,64742,0),
        (39407,47992,53462,57336,60312,62721,64742,0),
        (39409,47993,53463,57337,60313,62721,64743,0),
        (39412,47996,53464,57338,60313,62722,64743,0),
        (39415,47997,53465,57339,60314,62723,64744,0),
        (39417,47998,53466,57340,60315,62723,64744,0),
        (39419,48001,53468,57340,60315,62724,64745,0),
        (39423,48002,53469,57341,60316,62724,64745,0),
        (39425,48003,53470,57342,60317,62725,64746,0),
        (39427,48005,53471,57343,60317,62725,64746,0),
        (39431,48007,53472,57344,60318,62726,64746,0),
        (39433,48008,53473,57344,60318,62726,64747,0),
        (39435,48010,53474,57345,60319,62727,64747,0),
        (39438,48012,53475,57346,60320,62727,64748,0),
        (39441,48013,53476,57347,60320,62728,64748,0),
        (39444,48015,53477,57348,60321,62728,64749,0),
        (39446,48016,53479,57349,60322,62729,64749,0),
        (39449,48018,53480,57349,60322,62729,64750,0),
        (39452,48020,53481,57350,60323,62730,64750,0),
        (39454,48021,53482,57351,60324,62731,64751,0),
        (39456,48023,53483,57352,60324,62731,64751,0),
        (39460,48025,53484,57353,60325,62732,64752,0),
        (39462,48026,53485,57353,60326,62732,64752,0),
        (39464,48028,53486,57354,60326,62733,64752,0),
        (39468,48030,53487,57355,60327,62733,64753,0),
        (39470,48031,53488,57356,60327,62734,64753,0),
        (39472,48033,53489,57357,60328,62734,64754,0),
        (39475,48035,53491,57358,60329,62735,64754,0),
        (39478,48036,53492,57358,60329,62735,64755,0),
        (39480,48038,53493,57359,60330,62736,64755,0),
        (39483,48039,53494,57360,60331,62736,64756,0),
        (39486,48041,53495,57361,60331,62737,64756,0),
        (39488,48043,53496,57362,60332,62738,64757,0),
        (39491,48044,53497,57363,60333,62738,64757,0),
        (39493,48046,53498,57363,60333,62739,64757,0),
        (39496,48048,53499,57364,60334,62739,64758,0),
        (39499,48049,53500,57365,60335,62740,64758,0),
        (39501,48050,53502,57366,60335,62740,64759,0),
        (39505,48053,53503,57367,60336,62741,64759,0),
        (39507,48054,53504,57367,60336,62741,64760,0),
        (39509,48055,53505,57368,60337,62742,64760,0),
        (39511,48058,53506,57369,60338,62742,64760,0),
        (39515,48059,53507,57370,60338,62743,64761,0),
        (39517,48060,53508,57370,60339,62743,64761,0),
        (39519,48062,53510,57372,60340,62744,64762,0),
        (39523,48064,53510,57372,60340,62744,64762,0),
        (39525,48065,53511,57373,60341,62745,64763,0),
        (39528,48067,53512,57374,60342,62746,64763,0),
        (39530,48069,53514,57375,60342,62746,64764,0),
        (39533,48070,53515,57375,60343,62746,64764,0),
        (39536,48072,53516,57376,60344,62747,64765,0),
        (39538,48073,53517,57377,60344,62748,64765,0),
        (39541,48075,53518,57378,60345,62748,64765,0),
        (39544,48077,53519,57379,60345,62749,64766,0),
        (39546,48078,53520,57380,60346,62749,64766,0),
        (39548,48080,53522,57380,60347,62750,64767,0),
        (39552,48082,53522,57381,60347,62750,64767,0),
        (39554,48083,53523,57382,60348,62751,64768,0),
        (39556,48084,53525,57383,60349,62751,64768,0),
        (39560,48087,53526,57384,60349,62752,64769,0),
        (39562,48088,53527,57384,60350,62753,64769,0),
        (39564,48089,53528,57385,60351,62753,64770,0),
        (39567,48092,53529,57386,60351,62753,64770,0),
        (39570,48093,53530,57387,60352,62754,64771,0),
        (39572,48094,53531,57388,60353,62755,64771,0),
        (39575,48096,53533,57389,60353,62755,64771,0),
        (39578,48098,53533,57389,60354,62756,64772,0),
        (39580,48099,53534,57390,60354,62756,64772,0),
        (39583,48101,53535,57391,60355,62757,64773,0),
        (39585,48103,53537,57392,60356,62757,64773,0),
        (39588,48104,53538,57393,60356,62758,64774,0),
        (39591,48106,53539,57393,60357,62758,64774,0),
        (39593,48107,53540,57394,60358,62759,64775,0),
        (39596,48109,53541,57395,60358,62759,64775,0),
        (39599,48111,53542,57396,60359,62760,64776,0),
        (39601,48112,53543,57397,60360,62761,64776,0),
        (39603,48114,53544,57398,60360,62761,64776,0),
        (39607,48116,53545,57398,60361,62761,64777,0),
        (39609,48117,53546,57399,60362,62762,64777,0),
        (39611,48119,53548,57400,60362,62763,64778,0),
        (39615,48121,53549,57401,60363,62763,64778,0),
        (39617,48122,53550,57401,60364,62764,64779,0),
        (39619,48123,53551,57403,60364,62764,64779,0),
        (39622,48126,53552,57403,60365,62765,64780,0),
        (39625,48127,53553,57404,60365,62765,64780,0),
        (39627,48128,53554,57405,60366,62766,64781,0),
        (39630,48130,53555,57406,60367,62766,64781,0),
        (39633,48132,53556,57406,60367,62767,64781,0),
        (39635,48133,53557,57407,60368,62768,64782,0),
        (39638,48135,53558,57408,60369,62768,64782,0),
        (39640,48137,53560,57409,60369,62768,64783,0),
        (39643,48138,53561,57410,60370,62769,64783,0),
        (39646,48140,53562,57410,60371,62770,64784,0),
        (39648,48141,53563,57411,60371,62770,64784,0),
        (39651,48143,53564,57412,60372,62771,64785,0),
        (39654,48145,53565,57413,60373,62771,64785,0),
        (39656,48146,53566,57414,60373,62772,64786,0),
        (39658,48148,53567,57415,60374,62772,64786,0),
        (39662,48150,53568,57415,60375,62773,64787,0),
        (39664,48151,53569,57416,60375,62773,64787,0),
        (39666,48152,53571,57417,60376,62774,64787,0),
        (39670,48155,53572,57418,60376,62774,64788,0),
        (39672,48156,53573,57419,60377,62775,64788,0),
        (39674,48157,53574,57420,60378,62775,64789,0),
        (39676,48159,53575,57420,60378,62776,64789,0),
        (39680,48161,53576,57421,60379,62776,64790,0),
        (39682,48162,53577,57422,60380,62777,64790,0),
        (39684,48164,53578,57423,60380,62778,64791,0),
        (39688,48166,53579,57424,60381,62778,64791,0),
        (39690,48167,53580,57424,60382,62779,64792,0),
        (39692,48169,53581,57425,60382,62779,64792,0),
        (39695,48171,53583,57426,60383,62780,64792,0),
        (39698,48172,53584,57427,60384,62780,64793,0),
        (39700,48174,53585,57427,60384,62781,64793,0),
        (39703,48175,53586,57429,60385,62781,64794,0),
        (39706,48177,53587,57429,60386,62782,64794,0),
        (39708,48179,53588,57430,60386,62782,64795,0),
        (39711,48180,53589,57431,60387,62783,64795,0),
        (39713,48182,53590,57432,60387,62783,64795,0),
        (39716,48183,53591,57432,60388,62784,64796,0),
        (39719,48185,53592,57433,60389,62785,64796,0),
        (39721,48186,53594,57434,60389,62785,64797,0),
        (39724,48188,53595,57435,60390,62785,64797,0),
        (39727,48190,53596,57436,60391,62786,64798,0),
        (39729,48191,53597,57437,60391,62787,64798,0),
        (39731,48193,53598,57437,60392,62787,64799,0),
        (39735,48195,53599,57438,60393,62788,64799,0),
        (39737,48196,53600,57439,60393,62788,64800,0),
        (39739,48198,53601,57440,60394,62789,64800,0),
        (39742,48200,53602,57441,60395,62789,64800,0),
        (39745,48201,53603,57441,60395,62790,64801,0),
        (39747,48202,53604,57442,60396,62790,64801,0),
        (39749,48205,53606,57443,60397,62791,64802,0),
        (39753,48206,53607,57444,60397,62791,64802,0),
        (39755,48207,53607,57444,60398,62792,64803,0),
        (39757,48209,53609,57446,60398,62792,64803,0),
        (39761,48211,53610,57446,60399,62793,64804,0),
        (39763,48212,53611,57447,60400,62794,64804,0),
        (39765,48214,53612,57448,60400,62794,64805,0),
        (39768,48216,53613,57449,60401,62795,64805,0),
        (39771,48217,53614,57449,60402,62795,64806,0),
        (39773,48219,53615,57450,60402,62796,64806,0),
        (39775,48220,53617,57451,60403,62796,64806,0),
        (39779,48222,53617,57452,60404,62797,64807,0),
        (39781,48224,53618,57453,60404,62797,64807,0),
        (39783,48225,53619,57454,60405,62798,64808,0),
        (39786,48227,53621,57454,60406,62798,64808,0),
        (39789,48228,53622,57455,60406,62799,64809,0),
        (39791,48230,53623,57456,60407,62799,64809,0),
        (39794,48231,53624,57457,60407,62800,64810,0),
        (39797,48233,53625,57458,60408,62800,64810,0),
        (39799,48235,53626,57458,60409,62801,64811,0),
        (39802,48236,53627,57459,60409,62802,64811,0),
        (39804,48238,53628,57460,60410,62802,64811,0),
        (39807,48240,53629,57461,60411,62802,64812,0),
        (39810,48241,53630,57462,60411,62803,64812,0),
        (39812,48243,53632,57463,60412,62804,64813,0),
        (39815,48245,53633,57463,60413,62804,64813,0),
        (39818,48246,53634,57464,60413,62805,64814,0),
        (39820,48247,53635,57465,60414,62805,64814,0),
        (39823,48250,53636,57466,60415,62806,64815,0),
        (39825,48251,53637,57466,60415,62806,64815,0),
        (39828,48252,53638,57468,60416,62807,64816,0),
        (39830,48254,53639,57468,60416,62807,64816,0),
        (39833,48256,53640,57469,60417,62808,64817,0),
        (39836,48257,53641,57470,60418,62809,64817,0),
        (39838,48259,53643,57471,60418,62809,64817,0),
        (39841,48261,53644,57471,60419,62809,64818,0),
        (39844,48262,53645,57472,60420,62810,64818,0),
        (39846,48264,53646,57473,60420,62811,64819,0),
        (39848,48266,53647,57474,60421,62811,64819,0),
        (39852,48267,53648,57475,60422,62812,64820,0),
        (39854,48268,53649,57475,60422,62812,64820,0),
        (39856,48270,53650,57476,60423,62813,64820,0),
        (39859,48272,53651,57477,60424,62813,64821,0),
        (39862,48273,53652,57478,60424,62814,64821,0),
        (39864,48275,53653,57479,60425,62814,64822,0),
        (39866,48277,53655,57480,60425,62815,64822,0),
        (39870,48278,53655,57480,60426,62815,64823,0),
        (39872,48280,53656,57481,60427,62816,64823,0),
        (39874,48281,53658,57482,60427,62816,64824,0),
        (39878,48283,53659,57483,60428,62817,64824,0),
        (39880,48285,53660,57483,60429,62818,64825,0),
        (39882,48286,53661,57485,60429,62818,64825,0),
        (39884,48288,53662,57485,60430,62819,64825,0),
        (39888,48289,53663,57486,60431,62819,64826,0),
        (39890,48291,53664,57487,60431,62820,64826,0),
        (39892,48292,53665,57488,60432,62820,64827,0),
        (39896,48294,53666,57488,60432,62821,64827,0),
        (39898,48296,53667,57489,60433,62821,64828,0),
        (39900,48297,53668,57490,60434,62822,64828,0),
        (39902,48299,53670,57491,60434,62822,64829,0),
        (39906,48301,53671,57492,60435,62823,64829,0),
        (39908,48302,53672,57492,60436,62823,64830,0),
        (39910,48303,53673,57493,60436,62824,64830,0),
        (39914,48306,53674,57494,60437,62824,64830,0),
        (39916,48307,53675,57495,60438,62825,64831,0),
        (39918,48308,53676,57496,60438,62825,64831,0),
        (39921,48310,53677,57497,60439,62826,64832,0),
        (39924,48312,53678,57497,60440,62826,64832,0),
        (39926,48313,53679,57498,60440,62827,64833,0),
        (39928,48315,53681,57499,60441,62828,64833,0),
        (39932,48317,53682,57500,60441,62828,64834,0),
        (39934,48318,53682,57500,60442,62829,64834,0),
        (39936,48320,53683,57501,60443,62829,64835,0),
        (39939,48322,53685,57502,60443,62830,64835,0),
        (39942,48323,53686,57503,60444,62830,64836,0),
        (39944,48324,53687,57504,60445,62831,64836,0),
        (39947,48326,53688,57505,60445,62831,64836,0),
        (39950,48328,53689,57505,60446,62832,64837,0),
        (39952,48329,53690,57506,60447,62832,64837,0),
        (39954,48331,53691,57507,60447,62833,64838,0),
        (39957,48333,53692,57508,60448,62833,64838,0),
        (39960,48334,53693,57509,60448,62834,64839,0),
        (39962,48336,53694,57509,60449,62835,64839,0),
        (39965,48337,53696,57510,60450,62835,64840,0),
        (39968,48339,53697,57511,60450,62835,64840,0),
        (39970,48340,53698,57512,60451,62836,64840,0),
        (39973,48342,53699,57513,60452,62837,64841,0),
        (39975,48344,53700,57513,60452,62837,64841,0),
        (39978,48345,53701,57514,60453,62838,64842,0),
        (39980,48347,53702,57515,60454,62838,64842,0),
        (39983,48348,53703,57516,60454,62839,64843,0),
        (39986,48350,53704,57517,60455,62839,64843,0),
        (39988,48352,53705,57517,60455,62840,64844,0),
        (39991,48353,53706,57518,60456,62840,64844,0),
        (39993,48355,53708,57519,60457,62841,64844,0),
        (39996,48356,53709,57520,60457,62841,64845,0),
        (39998,48358,53709,57521,60458,62842,64845,0),
        (40001,48359,53711,57522,60459,62842,64846,0),
        (40004,48361,53712,57522,60459,62843,64846,0),
        (40006,48363,53713,57523,60460,62844,64847,0),
        (40009,48364,53714,57524,60461,62844,64847,0),
        (40011,48366,53715,57525,60461,62845,64848,0),
        (40014,48368,53716,57525,60462,62845,64848,0),
        (40016,48369,53717,57526,60463,62846,64849,0),
        (40019,48370,53718,57527,60463,62846,64849,0),
        (40022,48372,53719,57528,60464,62847,64849,0),
        (40024,48374,53720,57529,60464,62847,64850,0),
        (40027,48375,53721,57530,60465,62848,64850,0),
        (40029,48377,53723,57530,60466,62848,64851,0),
        (40032,48379,53724,57531,60466,62849,64851,0),
        (40034,48380,53725,57532,60467,62849,64852,0),
        (40037,48382,53726,57533,60468,62850,64852,0),
        (40040,48384,53727,57534,60468,62850,64853,0),
        (40042,48385,53728,57534,60469,62851,64853,0),
        (40045,48386,53729,57535,60470,62851,64854,0),
        (40047,48388,53730,57536,60470,62852,64854,0),
        (40050,48390,53731,57537,60471,62852,64855,0),
        (40052,48391,53732,57537,60472,62853,64855,0),
        (40055,48393,53734,57539,60472,62854,64855,0),
        (40058,48395,53734,57539,60473,62854,64856,0),
        (40060,48396,53735,57540,60473,62855,64856,0),
        (40063,48397,53736,57541,60474,62855,64857,0),
        (40065,48400,53738,57542,60475,62856,64857,0),
        (40068,48401,53739,57542,60475,62856,64858,0),
        (40070,48402,53740,57543,60476,62857,64858,0),
        (40073,48404,53741,57544,60477,62857,64858,0),
        (40076,48406,53742,57545,60477,62858,64859,0),
        (40078,48407,53743,57546,60478,62858,64859,0),
        (40081,48409,53744,57547,60479,62859,64860,0),
        (40083,48411,53745,57547,60479,62859,64860,0),
        (40086,48412,53746,57548,60480,62860,64861,0),
        (40088,48413,53747,57549,60481,62861,64861,0),
        (40091,48415,53749,57550,60481,62861,64862,0),
        (40094,48417,53750,57551,60482,62861,64862,0),
        (40096,48418,53750,57551,60482,62862,64863,0),
        (40098,48420,53751,57552,60483,62863,64863,0),
        (40101,48422,53753,57553,60484,62863,64863,0),
        (40104,48423,53754,57554,60484,62864,64864,0),
        (40106,48425,53755,57554,60485,62864,64864,0),
        (40109,48426,53756,57555,60486,62865,64865,0),
        (40112,48428,53757,57556,60486,62865,64865,0),
        (40114,48429,53758,57557,60487,62866,64866,0),
        (40116,48431,53759,57558,60488,62866,64866,0),
        (40119,48433,53760,57559,60488,62867,64867,0),
        (40122,48434,53761,57559,60489,62867,64867,0),
        (40124,48436,53762,57560,60490,62868,64868,0),
        (40127,48437,53764,57561,60490,62868,64868,0),
        (40130,48439,53765,57562,60491,62869,64868,0),
        (40132,48440,53766,57562,60491,62870,64869,0),
        (40134,48442,53766,57564,60492,62870,64869,0),
        (40137,48444,53768,57564,60493,62870,64870,0),
        (40140,48445,53769,57565,60493,62871,64870,0),
        (40142,48447,53770,57566,60494,62872,64871,0),
        (40144,48448,53771,57567,60495,62872,64871,0),
        (40148,48450,53772,57567,60495,62873,64872,0),
        (40150,48452,53773,57568,60496,62873,64872,0),
        (40152,48453,53774,57569,60497,62874,64873,0),
        (40154,48455,53775,57570,60497,62874,64873,0),
        (40158,48456,53776,57571,60498,62875,64873,0),
        (40160,48458,53777,57571,60499,62875,64874,0),
        (40162,48459,53779,57572,60499,62876,64874,0),
        (40166,48461,53780,57573,60500,62876,64875,0),
        (40168,48463,53781,57574,60500,62877,64875,0),
        (40170,48464,53782,57575,60501,62877,64876,0),
        (40172,48466,53783,57575,60502,62878,64876,0),
        (40176,48467,53784,57576,60502,62878,64877,0),
        (40178,48469,53785,57577,60503,62879,64877,0),
        (40180,48470,53786,57578,60504,62879,64877,0),
        (40184,48472,53787,57579,60504,62880,64878,0),
        (40186,48474,53788,57579,60505,62881,64878,0),
        (40188,48475,53789,57580,60506,62881,64879,0),
        (40190,48477,53790,57581,60506,62882,64879,0),
        (40194,48478,53791,57582,60507,62882,64880,0),
        (40196,48480,53792,57582,60508,62883,64880,0),
        (40198,48481,53794,57584,60508,62883,64881,0),
        (40201,48483,53795,57584,60509,62884,64881,0),
        (40204,48485,53796,57585,60509,62884,64882,0),
        (40206,48486,53797,57586,60510,62885,64882,0),
        (40208,48488,53798,57587,60511,62885,64882,0),
        (40211,48490,53799,57587,60511,62886,64883,0),
        (40214,48491,53800,57588,60512,62886,64883,0),
        (40216,48492,53801,57589,60513,62887,64884,0),
        (40219,48494,53802,57590,60513,62887,64884,0),
        (40222,48496,53803,57591,60514,62888,64885,0),
        (40224,48497,53804,57592,60514,62889,64885,0),
        (40226,48499,53805,57592,60515,62889,64886,0),
        (40229,48501,53806,57593,60516,62889,64886,0),
        (40232,48502,53807,57594,60516,62890,64887,0),
        (40234,48503,53809,57595,60517,62891,64887,0),
        (40237,48505,53810,57595,60518,62891,64887,0),
        (40239,48507,53811,57596,60518,62892,64888,0),
        (40242,48508,53812,57597,60519,62892,64888,0),
        (40244,48510,53813,57598,60520,62893,64889,0),
        (40247,48512,53814,57599,60520,62893,64889,0),
        (40249,48513,53815,57599,60521,62894,64890,0),
        (40252,48514,53816,57600,60521,62894,64890,0),
        (40255,48516,53817,57601,60522,62895,64890,0),
        (40257,48518,53818,57602,60523,62895,64891,0),
        (40259,48519,53819,57603,60523,62896,64891,0),
        (40262,48521,53820,57604,60524,62896,64892,0),
        (40265,48523,53821,57604,60525,62897,64892,0),
        (40267,48524,53822,57605,60525,62898,64893,0),
        (40269,48525,53824,57606,60526,62898,64893,0),
        (40273,48527,53825,57607,60526,62898,64894,0),
        (40275,48529,53826,57607,60527,62899,64894,0),
        (40277,48530,53827,57608,60528,62900,64895,0),
        (40279,48532,53828,57609,60528,62900,64895,0),
        (40283,48534,53829,57610,60529,62901,64896,0),
        (40285,48535,53830,57611,60530,62901,64896,0),
        (40287,48536,53831,57612,60530,62902,64896,0),
        (40291,48538,53832,57612,60531,62902,64897,0),
        (40293,48540,53833,57613,60531,62903,64897,0),
        (40295,48541,53834,57614,60532,62903,64898,0),
        (40297,48543,53835,57615,60533,62904,64898,0),
        (40301,48545,53836,57615,60533,62904,64899,0),
        (40303,48546,53837,57616,60534,62905,64899,0),
        (40305,48547,53839,57617,60535,62905,64900,0),
        (40308,48549,53840,57618,60535,62906,64900,0),
        (40311,48551,53841,57619,60536,62907,64901,0),
        (40313,48552,53842,57620,60537,62907,64901,0),
        (40315,48554,53843,57620,60537,62907,64901,0),
        (40318,48556,53844,57621,60538,62908,64902,0),
        (40321,48557,53845,57622,60539,62909,64902,0),
        (40323,48558,53846,57623,60539,62909,64903,0),
        (40326,48560,53847,57623,60540,62910,64903,0),
        (40328,48562,53848,57624,60540,62910,64904,0),
        (40331,48563,53849,57625,60541,62911,64904,0),
        (40333,48565,53850,57626,60542,62911,64904,0),
        (40336,48567,53851,57627,60542,62912,64905,0),
        (40338,48568,53852,57627,60543,62912,64905,0),
        (40341,48569,53854,57628,60544,62913,64906,0),
        (40344,48571,53855,57629,60544,62913,64906,0),
        (40346,48573,53856,57630,60545,62914,64907,0),
        (40348,48574,53857,57631,60546,62914,64907,0),
        (40351,48576,53858,57632,60546,62915,64908,0),
        (40354,48578,53859,57632,60547,62915,64908,0),
        (40356,48579,53860,57633,60548,62916,64909,0),
        (40358,48580,53861,57634,60548,62916,64909,0),
        (40362,48582,53862,57635,60549,62917,64909,0),
        (40364,48584,53863,57635,60549,62918,64910,0),
        (40366,48585,53864,57636,60550,62918,64910,0),
        (40368,48587,53865,57637,60551,62919,64911,0),
        (40372,48589,53866,57638,60551,62919,64911,0),
        (40374,48590,53867,57639,60552,62920,64912,0),
        (40376,48591,53869,57640,60553,62920,64912,0),
        (40379,48593,53870,57640,60553,62921,64913,0),
        (40382,48595,53871,57641,60554,62921,64913,0),
        (40384,48596,53871,57642,60555,62922,64913,0),
        (40386,48598,53873,57643,60555,62922,64914,0),
        (40389,48599,53874,57643,60556,62923,64914,0),
        (40392,48601,53875,57644,60557,62923,64915,0),
        (40394,48602,53876,57645,60557,62924,64915,0),
        (40397,48604,53877,57646,60558,62924,64916,0),
        (40399,48606,53878,57647,60558,62925,64916,0),
        (40402,48607,53879,57648,60559,62925,64917,0),
        (40404,48609,53880,57648,60560,62926,64917,0),
        (40407,48610,53881,57649,60560,62926,64918,0),
        (40409,48612,53882,57650,60561,62927,64918,0),
        (40412,48613,53884,57651,60562,62928,64918,0),
        (40415,48615,53885,57651,60562,62928,64919,0),
        (40417,48617,53885,57652,60563,62929,64919,0),
        (40419,48618,53886,57653,60563,62929,64920,0),
        (40421,48620,53888,57654,60564,62930,64920,0),
        (40425,48621,53889,57655,60565,62930,64921,0),
        (40427,48623,53890,57655,60565,62931,64921,0),
        (40429,48624,53891,57656,60566,62931,64922,0),
        (40433,48626,53892,57657,60567,62932,64922,0),
        (40435,48628,53893,57658,60567,62932,64923,0),
        (40437,48629,53894,57659,60568,62933,64923,0),
        (40439,48631,53895,57659,60568,62933,64923,0),
        (40442,48632,53896,57660,60569,62934,64924,0),
        (40445,48634,53897,57661,60570,62934,64924,0),
        (40447,48635,53898,57662,60570,62935,64925,0),
        (40450,48637,53899,57663,60571,62935,64925,0),
        (40452,48638,53900,57663,60572,62936,64926,0),
        (40455,48640,53901,57664,60572,62936,64926,0),
        (40457,48642,53903,57665,60573,62937,64926,0),
        (40460,48643,53904,57666,60573,62937,64927,0),
        (40462,48645,53905,57666,60574,62938,64927,0),
        (40465,48646,53906,57668,60575,62939,64928,0),
        (40468,48648,53907,57668,60575,62939,64928,0),
        (40470,48649,53908,57669,60576,62940,64929,0),
        (40472,48651,53909,57670,60577,62940,64929,0),
        (40475,48653,53910,57671,60577,62941,64930,0),
        (40478,48654,53911,57671,60578,62941,64930,0),
        (40480,48656,53912,57672,60579,62942,64931,0),
        (40482,48657,53913,57673,60579,62942,64931,0),
        (40486,48659,53914,57674,60580,62943,64931,0),
        (40488,48660,53915,57674,60580,62943,64932,0),
        (40490,48662,53916,57676,60581,62944,64932,0),
        (40492,48664,53918,57676,60582,62944,64933,0),
        (40495,48665,53919,57677,60582,62945,64933,0),
        (40498,48666,53919,57678,60583,62945,64934,0),
        (40500,48668,53921,57679,60584,62946,64934,0),
        (40503,48670,53922,57679,60584,62946,64935,0),
        (40505,48671,53923,57680,60585,62947,64935,0),
        (40508,48673,53924,57681,60586,62948,64936,0),
        (40510,48675,53925,57682,60586,62948,64936,0),
        (40513,48676,53926,57682,60587,62948,64936,0),
        (40515,48677,53927,57684,60588,62949,64937,0),
        (40517,48679,53928,57684,60588,62950,64937,0),
        (40521,48681,53929,57685,60589,62950,64938,0),
        (40523,48682,53930,57686,60590,62951,64938,0),
        (40525,48683,53932,57687,60590,62951,64939,0),
        (40529,48686,53932,57687,60591,62952,64939,0),
        (40531,48687,53933,57688,60591,62952,64940,0),
        (40533,48688,53934,57689,60592,62953,64940,0),
        (40535,48690,53936,57690,60593,62953,64940,0),
        (40538,48692,53937,57690,60593,62954,64941,0),
        (40541,48693,53938,57691,60594,62954,64941,0),
        (40543,48694,53939,57692,60595,62955,64942,0),
        (40546,48696,53940,57693,60595,62955,64942,0),
        (40548,48698,53941,57694,60596,62956,64943,0),
        (40551,48699,53942,57695,60597,62957,64943,0),
        (40553,48701,53943,57695,60597,62957,64944,0),
        (40556,48703,53944,57696,60598,62957,64944,0),
        (40558,48704,53945,57697,60598,62958,64945,0),
        (40560,48705,53946,57698,60599,62959,64945,0),
        (40564,48707,53947,57698,60600,62959,64945,0),
        (40566,48709,53948,57699,60600,62960,64946,0),
        (40568,48710,53949,57700,60601,62960,64946,0),
        (40570,48712,53951,57701,60601,62961,64947,0),
        (40574,48713,53951,57702,60602,62961,64947,0),
        (40576,48715,53952,57702,60603,62962,64948,0),
        (40578,48716,53954,57703,60603,62962,64948,0),
        (40581,48718,53955,57704,60604,62963,64948,0),
        (40583,48720,53956,57705,60605,62963,64949,0),
        (40586,48721,53957,57706,60605,62964,64949,0),
        (40588,48723,53958,57706,60606,62964,64950,0),
        (40591,48724,53959,57707,60606,62965,64950,0),
        (40593,48726,53960,57708,60607,62965,64951,0),
        (40596,48727,53961,57709,60608,62966,64951,0),
        (40599,48729,53962,57710,60608,62966,64952,0),
        (40601,48730,53963,57710,60609,62967,64952,0),
        (40603,48732,53964,57711,60610,62968,64953,0),
        (40605,48734,53965,57712,60610,62968,64953,0),
        (40609,48735,53966,57713,60611,62968,64954,0),
        (40611,48736,53967,57713,60612,62969,64954,0),
        (40613,48738,53969,57714,60612,62970,64954,0),
        (40616,48740,53970,57715,60613,62970,64955,0),
        (40619,48741,53970,57716,60613,62971,64955,0),
        (40621,48743,53971,57717,60614,62971,64956,0),
        (40623,48745,53973,57718,60615,62972,64956,0),
        (40626,48746,53974,57718,60615,62972,64957,0),
        (40628,48747,53975,57719,60616,62973,64957,0),
        (40631,48749,53976,57720,60617,62973,64957,0),
        (40634,48751,53977,57721,60617,62974,64958,0),
        (40636,48752,53978,57721,60618,62974,64958,0),
        (40638,48753,53979,57722,60619,62975,64959,0),
        (40640,48755,53980,57723,60619,62975,64959,0),
        (40644,48757,53981,57724,60620,62976,64960,0),
        (40646,48758,53982,57725,60621,62977,64960,0),
        (40648,48760,53983,57726,60621,62977,64961,0),
        (40651,48762,53984,57726,60622,62977,64961,0),
        (40654,48763,53985,57727,60622,62978,64962,0),
        (40656,48764,53986,57728,60623,62979,64962,0),
        (40658,48766,53988,57729,60624,62979,64962,0),
        (40661,48768,53989,57729,60624,62979,64963,0),
        (40663,48769,53989,57730,60625,62980,64963,0),
        (40666,48770,53991,57731,60626,62981,64964,0),
        (40669,48772,53992,57732,60626,62981,64964,0),
        (40671,48774,53993,57733,60627,62982,64965,0),
        (40673,48775,53994,57734,60628,62982,64965,0),
        (40676,48777,53995,57734,60628,62983,64966,0),
        (40679,48778,53996,57735,60629,62983,64966,0),
        (40681,48780,53997,57736,60629,62984,64966,0),
        (40683,48781,53998,57737,60630,62984,64967,0),
        (40686,48783,53999,57737,60631,62985,64967,0),
        (40689,48785,54000,57738,60631,62985,64968,0),
        (40691,48786,54001,57739,60632,62986,64968,0),
        (40693,48788,54002,57740,60632,62986,64969,0),
        (40696,48789,54003,57741,60633,62987,64969,0),
        (40698,48791,54004,57741,60634,62988,64970,0),
        (40701,48792,54006,57742,60634,62988,64970,0),
        (40704,48794,54007,57743,60635,62988,64970,0),
        (40706,48795,54008,57744,60636,62989,64971,0),
        (40708,48797,54008,57745,60636,62990,64971,0),
        (40710,48799,54010,57745,60637,62990,64972,0),
        (40714,48800,54011,57746,60637,62990,64972,0),
        (40716,48801,54012,57747,60638,62991,64973,0),
        (40718,48803,54013,57748,60639,62992,64973,0),
        (40721,48805,54014,57748,60639,62992,64974,0),
        (40724,48806,54015,57749,60640,62993,64974,0),
        (40726,48808,54016,57750,60641,62993,64975,0),
        (40728,48810,54017,57751,60641,62994,64975,0),
        (40731,48811,54018,57752,60642,62994,64976,0),
        (40733,48812,54019,57752,60643,62995,64976,0),
        (40736,48814,54020,57753,60643,62995,64976,0),
        (40739,48816,54021,57754,60644,62996,64977,0),
        (40741,48817,54022,57755,60644,62996,64977,0),
        (40743,48818,54023,57756,60645,62997,64978,0),
        (40745,48820,54025,57756,60646,62997,64978,0),
        (40749,48822,54026,57757,60646,62998,64979,0),
        (40751,48823,54026,57758,60647,62999,64979,0),
        (40753,48824,54028,57759,60648,62999,64979,0),
        (40756,48826,54029,57760,60648,62999,64980,0),
        (40758,48828,54030,57760,60649,63000,64980,0),
        (40761,48829,54031,57761,60650,63001,64981,0),
        (40763,48831,54032,57762,60650,63001,64981,0),
        (40766,48832,54033,57763,60651,63001,64982,0),
        (40768,48834,54034,57763,60652,63002,64982,0),
        (40770,48835,54035,57764,60652,63003,64983,0),
        (40774,48837,54036,57765,60653,63003,64983,0),
        (40776,48839,54037,57766,60653,63004,64984,0),
        (40778,48840,54038,57767,60654,63004,64984,0),
        (40780,48842,54039,57768,60655,63005,64984,0),
        (40783,48843,54040,57768,60655,63005,64985,0),
        (40786,48845,54041,57769,60656,63006,64985,0),
        (40788,48846,54043,57770,60657,63006,64986,0),
        (40791,48848,54043,57771,60657,63007,64986,0),
        (40793,48849,54044,57771,60658,63007,64987,0),
        (40795,48851,54045,57772,60658,63008,64987,0),
        (40798,48853,54047,57773,60659,63008,64987,0),
        (40801,48854,54048,57774,60660,63009,64988,0),
        (40803,48855,54049,57774,60660,63010,64988,0),
        (40805,48857,54050,57775,60661,63010,64989,0),
        (40809,48859,54051,57776,60661,63010,64989,0),
        (40811,48860,54052,57777,60662,63011,64990,0),
        (40813,48861,54053,57778,60663,63012,64990,0),
        (40815,48863,54054,57779,60663,63012,64991,0),
        (40818,48865,54055,57779,60664,63012,64991,0),
        (40820,48866,54056,57780,60665,63013,64992,0),
        (40823,48867,54057,57781,60665,63014,64992,0),
        (40826,48869,54058,57782,60666,63014,64992,0),
        (40828,48871,54059,57782,60666,63015,64993,0),
        (40830,48872,54060,57783,60667,63015,64993,0),
        (40832,48874,54061,57784,60668,63016,64994,0),
        (40836,48876,54062,57785,60668,63016,64994,0),
        (40838,48877,54063,57786,60669,63017,64995,0),
        (40840,48878,54065,57787,60670,63017,64995,0),
        (40843,48880,54066,57787,60670,63018,64995,0),
        (40845,48882,54067,57788,60671,63018,64996,0),
        (40848,48883,54067,57789,60672,63019,64996,0),
        (40850,48885,54069,57790,60672,63019,64997,0),
        (40853,48886,54070,57790,60673,63020,64997,0),
        (40855,48888,54071,57791,60674,63020,64998,0),
        (40857,48889,54072,57792,60674,63021,64998,0),
        (40861,48891,54073,57793,60675,63021,64999,0),
        (40863,48892,54074,57793,60675,63022,64999,0),
        (40865,48894,54075,57794,60676,63023,65000,0),
        (40867,48896,54076,57795,60677,63023,65000,0),
        (40870,48897,54077,57796,60677,63023,65001,0),
        (40873,48898,54078,57797,60678,63024,65001,0),
        (40875,48900,54079,57798,60679,63025,65001,0),
        (40878,48902,54080,57798,60679,63025,65002,0),
        (40880,48903,54081,57799,60680,63026,65002,0),
        (40882,48904,54082,57800,60680,63026,65003,0),
        (40884,48906,54084,57801,60681,63027,65003,0),
        (40888,48908,54084,57801,60682,63027,65004,0),
        (40890,48909,54085,57802,60682,63028,65004,0),
        (40892,48910,54087,57803,60683,63028,65004,0),
        (40895,48912,54088,57804,60684,63029,65005,0),
        (40897,48914,54089,57805,60684,63029,65005,0),
        (40900,48915,54089,57806,60685,63030,65006,0),
        (40902,48917,54091,57806,60685,63030,65006,0),
        (40905,48918,54092,57807,60686,63031,65007,0),
        (40907,48920,54093,57808,60687,63031,65007,0),
        (40909,48921,54094,57809,60687,63032,65008,0),
        (40913,48923,54095,57809,60688,63032,65008,0),
        (40915,48924,54096,57810,60688,63033,65009,0),
        (40917,48926,54097,57811,60689,63034,65009,0),
        (40919,48928,54098,57812,60690,63034,65009,0),
        (40922,48929,54099,57812,60690,63034,65010,0),
        (40924,48930,54100,57813,60691,63035,65010,0),
        (40927,48932,54101,57814,60692,63036,65011,0),
        (40930,48934,54102,57815,60692,63036,65011,0),
        (40932,48935,54103,57816,60693,63037,65012,0),
        (40934,48937,54104,57817,60694,63037,65012,0),
        (40936,48939,54106,57817,60694,63038,65012,0),
        (40940,48940,54106,57818,60695,63038,65013,0),
        (40942,48941,54107,57819,60696,63039,65013,0),
        (40944,48943,54109,57820,60696,63039,65014,0),
        (40947,48945,54110,57820,60697,63040,65014,0),
        (40949,48946,54111,57821,60697,63040,65015,0),
        (40951,48947,54111,57822,60698,63041,65015,0),
        (40954,48949,54113,57823,60699,63041,65016,0),
        (40957,48951,54114,57823,60699,63042,65016,0),
        (40959,48952,54115,57824,60700,63042,65017,0),
        (40961,48953,54116,57825,60701,63043,65017,0),
        (40964,48955,54117,57826,60701,63043,65017,0),
        (40967,48957,54118,57827,60702,63044,65018,0),
        (40969,48958,54119,57828,60702,63044,65018,0),
        (40971,48960,54120,57828,60703,63045,65019,0),
        (40974,48961,54121,57829,60704,63045,65019,0),
        (40976,48963,54122,57830,60704,63046,65020,0),
        (40978,48964,54123,57831,60705,63047,65020,0),
        (40982,48966,54124,57831,60706,63047,65020,0),
        (40984,48967,54125,57832,60706,63048,65021,0),
        (40986,48969,54126,57833,60707,63048,65021,0),
        (40988,48971,54128,57834,60707,63049,65022,0),
        (40991,48972,54128,57834,60708,63049,65022,0),
        (40994,48973,54129,57835,60709,63050,65023,0),
        (40996,48975,54131,57836,60709,63050,65023,0),
        (40999,48977,54132,57837,60710,63051,65024,0),
        (41001,48978,54133,57838,60710,63051,65024,0),
        (41003,48979,54133,57839,60711,63052,65025,0),
        (41005,48981,54135,57839,60712,63052,65025,0),
        (41009,48983,54136,57840,60712,63053,65026,0),
        (41011,48984,54137,57841,60713,63053,65026,0),
        (41013,48985,54138,57842,60714,63054,65026,0),
        (41016,48987,54139,57842,60714,63054,65027,0),
        (41018,48989,54140,57843,60715,63055,65027,0),
        (41020,48990,54141,57844,60716,63055,65028,0),
        (41023,48992,54142,57845,60716,63056,65028,0),
        (41026,48993,54143,57845,60717,63056,65029,0),
        (41028,48995,54144,57846,60718,63057,65029,0),
        (41030,48996,54145,57847,60718,63057,65029,0),
        (41033,48998,54146,57848,60719,63058,65030,0),
        (41036,48999,54147,57849,60719,63059,65030,0),
        (41038,49001,54148,57850,60720,63059,65031,0),
        (41040,49003,54149,57850,60721,63060,65031,0),
        (41043,49004,54150,57851,60721,63060,65032,0),
        (41045,49005,54151,57852,60722,63061,65032,0),
        (41047,49007,54153,57853,60723,63061,65033,0),
        (41051,49009,54154,57853,60723,63062,65033,0),
        (41053,49010,54155,57854,60724,63062,65034,0),
        (41055,49011,54155,57855,60724,63063,65034,0),
        (41057,49013,54157,57856,60725,63063,65034,0),
        (41060,49015,54158,57856,60726,63064,65035,0),
        (41062,49016,54159,57857,60726,63064,65035,0),
        (41065,49017,54160,57858,60727,63065,65036,0),
        (41068,49019,54161,57859,60727,63065,65036,0),
        (41070,49021,54162,57860,60728,63066,65037,0),
        (41072,49022,54163,57861,60729,63066,65037,0),
        (41074,49024,54164,57861,60729,63067,65037,0),
        (41077,49025,54165,57862,60730,63067,65038,0),
        (41080,49027,54166,57863,60731,63068,65038,0),
        (41082,49028,54167,57864,60731,63068,65039,0),
        (41085,49030,54168,57864,60732,63069,65039,0),
        (41087,49031,54169,57865,60732,63070,65040,0),
        (41089,49033,54170,57866,60733,63070,65040,0),
        (41091,49035,54171,57867,60734,63070,65041,0),
        (41095,49036,54172,57867,60734,63071,65041,0),
        (41097,49037,54173,57868,60735,63072,65041,0),
        (41099,49038,54175,57869,60736,63072,65042,0),
        (41102,49040,54176,57870,60736,63073,65042,0),
        (41104,49042,54176,57871,60737,63073,65043,0),
        (41106,49043,54177,57872,60738,63074,65043,0),
        (41109,49045,54179,57872,60738,63074,65044,0),
        (41112,49046,54180,57873,60739,63075,65044,0),
        (41114,49048,54181,57874,60740,63075,65045,0),
        (41116,49049,54182,57875,60740,63076,65045,0),
        (41119,49051,54183,57875,60741,63076,65045,0),
        (41121,49052,54184,57876,60741,63077,65046,0),
        (41124,49054,54185,57877,60742,63077,65046,0),
        (41126,49056,54186,57878,60743,63078,65047,0),
        (41129,49057,54187,57878,60743,63078,65047,0),
        (41131,49058,54188,57879,60744,63079,65048,0),
        (41133,49060,54189,57880,60744,63079,65048,0),
        (41136,49062,54190,57881,60745,63080,65049,0),
        (41139,49063,54191,57882,60746,63081,65049,0),
        (41141,49064,54192,57883,60746,63081,65049,0),
        (41143,49066,54193,57883,60747,63081,65050,0),
        (41146,49068,54194,57884,60747,63082,65050,0),
        (41148,49069,54195,57885,60748,63083,65051,0),
        (41150,49070,54196,57886,60749,63083,65051,0),
        (41153,49072,54197,57886,60749,63083,65052,0),
        (41156,49074,54198,57887,60750,63084,65052,0),
        (41158,49075,54199,57888,60751,63085,65053,0),
        (41160,49077,54201,57889,60751,63085,65053,0),
        (41163,49078,54201,57889,60752,63086,65054,0),
        (41165,49080,54202,57890,60753,63086,65054,0),
        (41167,49081,54204,57891,60753,63087,65054,0),
        (41171,49083,54205,57892,60754,63087,65055,0),
        (41173,49084,54206,57893,60754,63088,65055,0),
        (41175,49086,54206,57894,60755,63088,65056,0),
        (41177,49088,54208,57894,60756,63089,65056,0),
        (41180,49089,54209,57895,60756,63089,65057,0),
        (41182,49090,54210,57896,60757,63090,65057,0),
        (41184,49092,54211,57897,60758,63090,65057,0),
        (41188,49094,54212,57897,60758,63091,65058,0),
        (41190,49095,54213,57898,60759,63091,65058,0),
        (41192,49096,54214,57899,60760,63092,65059,0),
        (41195,49098,54215,57900,60760,63092,65059,0),
        (41197,49099,54216,57900,60761,63093,65060,0),
        (41199,49101,54217,57901,60761,63093,65060,0),
        (41202,49103,54218,57902,60762,63094,65061,0),
        (41205,49104,54219,57903,60763,63094,65061,0),
        (41207,49105,54220,57903,60763,63095,65062,0),
        (41209,49107,54221,57905,60764,63096,65062,0),
        (41212,49109,54222,57905,60764,63096,65062,0),
        (41214,49110,54223,57906,60765,63097,65063,0),
        (41216,49111,54224,57907,60766,63097,65063,0),
        (41219,49113,54226,57908,60766,63098,65064,0),
        (41222,49115,54226,57908,60767,63098,65064,0),
        (41224,49116,54227,57909,60768,63099,65065,0),
        (41226,49117,54229,57910,60768,63099,65065,0),
        (41229,49119,54230,57911,60769,63100,65065,0),
        (41231,49121,54231,57911,60769,63100,65066,0),
        (41234,49122,54231,57912,60770,63101,65066,0),
        (41236,49124,54233,57913,60771,63101,65067,0),
        (41239,49125,54234,57914,60771,63102,65067,0),
        (41241,49127,54235,57914,60772,63102,65068,0),
        (41243,49128,54236,57915,60773,63103,65068,0),
        (41246,49130,54237,57916,60773,63103,65069,0),
        (41248,49131,54238,57917,60774,63104,65069,0),
        (41251,49132,54239,57918,60775,63104,65070,0),
        (41253,49134,54240,57919,60775,63105,65070,0),
        (41256,49136,54241,57919,60776,63105,65070,0),
        (41258,49137,54242,57920,60776,63106,65071,0),
        (41260,49138,54243,57921,60777,63106,65071,0),
        (41263,49140,54244,57922,60778,63107,65072,0),
        (41265,49142,54245,57922,60778,63108,65072,0),
        (41268,49143,54246,57923,60779,63108,65073,0),
        (41270,49145,54247,57924,60779,63108,65073,0),
        (41273,49146,54248,57925,60780,63109,65074,0),
        (41275,49148,54249,57925,60781,63110,65074,0),
        (41277,49149,54251,57926,60781,63110,65074,0),
        (41280,49151,54251,57927,60782,63111,65075,0),
        (41282,49152,54252,57928,60782,63111,65075,0),
        (41285,49154,54253,57929,60783,63112,65076,0),
        (41287,49156,54255,57929,60784,63112,65076,0),
        (41290,49157,54256,57930,60784,63113,65077,0),
        (41292,49158,54256,57931,60785,63113,65077,0),
        (41294,49160,54258,57932,60786,63114,65077,0),
        (41297,49161,54259,57933,60786,63114,65078,0),
        (41299,49163,54260,57933,60787,63115,65078,0),
        (41302,49164,54261,57934,60788,63115,65079,0),
        (41304,49166,54262,57935,60788,63116,65079,0),
        (41307,49167,54263,57936,60789,63116,65080,0),
        (41309,49169,54264,57936,60790,63117,65080,0),
        (41311,49170,54265,57937,60790,63117,65081,0),
        (41314,49172,54266,57938,60791,63118,65081,0),
        (41316,49173,54267,57939,60791,63118,65082,0),
        (41319,49175,54268,57940,60792,63119,65082,0),
        (41321,49177,54269,57940,60793,63119,65082,0),
        (41324,49178,54270,57941,60793,63120,65083,0),
        (41326,49179,54271,57942,60794,63121,65083,0),
        (41328,49181,54272,57943,60795,63121,65084,0),
        (41331,49183,54273,57943,60795,63121,65084,0),
        (41333,49184,54274,57944,60796,63122,65085,0),
        (41336,49185,54275,57945,60796,63123,65085,0),
        (41338,49187,54276,57946,60797,63123,65085,0),
        (41341,49188,54277,57947,60798,63123,65086,0),
        (41343,49190,54278,57947,60798,63124,65086,0),
        (41345,49191,54280,57948,60799,63125,65087,0),
        (41348,49193,54280,57949,60799,63125,65087,0),
        (41350,49194,54281,57950,60800,63126,65088,0),
        (41353,49196,54282,57951,60801,63126,65088,0),
        (41355,49198,54284,57951,60801,63127,65089,0),
        (41358,49199,54285,57952,60802,63127,65089,0),
        (41360,49200,54285,57953,60803,63128,65089,0),
        (41362,49202,54287,57954,60803,63128,65090,0),
        (41365,49204,54288,57954,60804,63129,65090,0),
        (41367,49205,54289,57955,60804,63129,65091,0),
        (41369,49206,54289,57956,60805,63130,65091,0),
        (41372,49208,54291,57957,60806,63130,65092,0),
        (41375,49209,54292,57957,60806,63131,65092,0),
        (41377,49211,54293,57958,60807,63131,65093,0),
        (41379,49212,54294,57959,60808,63132,65093,0),
        (41382,49214,54295,57960,60808,63132,65093,0),
        (41384,49215,54296,57961,60809,63133,65094,0),
        (41386,49217,54297,57962,60810,63133,65094,0),
        (41388,49219,54298,57962,60810,63134,65095,0),
        (41392,49220,54299,57963,60811,63134,65095,0),
        (41394,49221,54300,57964,60811,63135,65096,0),
        (41396,49223,54301,57965,60812,63135,65096,0),
        (41399,49225,54302,57965,60813,63136,65096,0),
        (41401,49226,54303,57966,60813,63137,65097,0),
        (41403,49227,54304,57967,60814,63137,65097,0),
        (41405,49229,54305,57968,60814,63138,65098,0),
        (41409,49230,54306,57968,60815,63138,65098,0),
        (41411,49232,54307,57969,60816,63139,65099,0),
        (41413,49233,54308,57970,60816,63139,65099,0),
        (41416,49235,54309,57971,60817,63140,65100,0),
        (41418,49236,54310,57971,60817,63140,65100,0),
        (41420,49238,54311,57972,60818,63141,65101,0),
        (41422,49240,54313,57973,60819,63141,65101,0),
        (41425,49241,54313,57974,60819,63142,65102,0),
        (41428,49242,54314,57975,60820,63142,65102,0),
        (41430,49244,54316,57976,60821,63143,65102,0),
        (41433,49246,54317,57976,60821,63143,65103,0),
        (41435,49247,54318,57977,60822,63144,65103,0),
        (41437,49248,54318,57978,60823,63144,65104,0),
        (41439,49250,54320,57979,60823,63145,65104,0),
        (41442,49251,54321,57979,60824,63145,65105,0),
        (41444,49253,54322,57980,60824,63146,65105,0),
        (41447,49254,54323,57981,60825,63146,65105,0),
        (41450,49256,54324,57982,60826,63147,65106,0),
        (41452,49257,54325,57982,60826,63147,65106,0),
        (41454,49259,54326,57983,60827,63148,65107,0),
        (41456,49261,54327,57984,60827,63148,65107,0),
        (41459,49262,54328,57985,60828,63149,65108,0),
        (41461,49263,54329,57985,60829,63150,65108,0),
        (41463,49264,54330,57986,60829,63150,65108,0),
        (41467,49266,54331,57987,60830,63150,65109,0),
        (41469,49268,54332,57988,60830,63151,65109,0),
        (41471,49269,54333,57989,60831,63152,65110,0),
        (41473,49271,54334,57989,60832,63152,65110,0),
        (41476,49272,54335,57990,60832,63152,65111,0),
        (41478,49274,54336,57991,60833,63153,65111,0),
        (41480,49275,54337,57992,60834,63154,65112,0),
        (41483,49277,54338,57993,60834,63154,65112,0),
        (41486,49278,54339,57993,60835,63155,65113,0),
        (41488,49280,54340,57994,60836,63155,65113,0),
        (41490,49281,54341,57995,60836,63156,65113,0),
        (41493,49283,54342,57996,60837,63156,65114,0),
        (41495,49284,54343,57996,60838,63157,65114,0),
        (41497,49285,54345,57997,60838,63157,65115,0),
        (41500,49287,54345,57998,60839,63158,65115,0),
        (41502,49289,54346,57999,60839,63158,65116,0),
        (41504,49290,54347,58000,60840,63159,65116,0),
        (41507,49292,54349,58000,60841,63159,65116,0),
        (41510,49293,54350,58001,60841,63160,65117,0),
        (41512,49295,54350,58002,60842,63160,65117,0),
        (41514,49296,54352,58003,60842,63161,65118,0),
        (41517,49298,54353,58003,60843,63161,65118,0),
        (41519,49299,54354,58004,60844,63162,65119,0),
        (41521,49300,54354,58005,60844,63162,65119,0),
        (41523,49302,54356,58006,60845,63163,65120,0),
        (41527,49304,54357,58006,60845,63163,65120,0),
        (41529,49305,54358,58007,60846,63164,65120,0),
        (41531,49306,54359,58008,60847,63164,65121,0),
        (41534,49308,54360,58009,60847,63165,65121,0),
        (41536,49310,54361,58010,60848,63166,65122,0),
        (41538,49311,54362,58011,60849,63166,65122,0),
        (41540,49313,54363,58011,60849,63166,65123,0),
        (41543,49314,54364,58012,60850,63167,65123,0),
        (41545,49315,54365,58013,60851,63168,65124,0),
        (41548,49317,54366,58014,60851,63168,65124,0),
        (41551,49319,54367,58014,60852,63169,65124,0),
        (41553,49320,54368,58015,60852,63169,65125,0),
        (41555,49321,54369,58016,60853,63170,65125,0),
        (41557,49323,54370,58017,60854,63170,65126,0),
        (41560,49325,54371,58017,60854,63171,65126,0),
        (41562,49326,54372,58018,60855,63171,65127,0),
        (41564,49327,54373,58019,60855,63172,65127,0),
        (41567,49329,54374,58020,60856,63172,65127,0),
        (41570,49330,54375,58020,60857,63173,65128,0),
        (41572,49332,54376,58021,60857,63173,65128,0),
        (41574,49334,54377,58022,60858,63174,65129,0),
        (41577,49335,54378,58023,60858,63174,65129,0),
        (41579,49336,54379,58023,60859,63175,65130,0),
        (41581,49338,54381,58024,60860,63175,65130,0),
        (41584,49339,54381,58025,60860,63176,65131,0),
        (41586,49341,54382,58026,60861,63176,65131,0),
        (41588,49342,54383,58027,60862,63177,65132,0),
        (41591,49344,54385,58028,60862,63177,65132,0),
        (41594,49345,54385,58028,60863,63178,65132,0),
        (41596,49347,54386,58029,60864,63178,65133,0),
        (41598,49348,54388,58030,60864,63179,65133,0),
        (41601,49350,54389,58031,60865,63179,65134,0),
        (41603,49351,54390,58031,60865,63180,65134,0),
        (41605,49352,54390,58032,60866,63181,65135,0),
        (41607,49354,54392,58033,60867,63181,65135,0),
        (41610,49356,54393,58034,60867,63181,65136,0),
        (41612,49357,54394,58034,60868,63182,65136,0),
        (41615,49358,54395,58035,60869,63183,65136,0),
        (41618,49360,54396,58036,60869,63183,65137,0),
        (41620,49362,54397,58037,60870,63184,65137,0),
        (41622,49363,54398,58038,60870,63184,65138,0),
        (41624,49365,54399,58038,60871,63185,65138,0),
        (41627,49366,54400,58039,60871,63185,65139,0),
        (41629,49367,54401,58040,60872,63186,65139,0),
        (41631,49369,54402,58041,60873,63186,65139,0),
        (41634,49371,54403,58041,60873,63187,65140,0),
        (41637,49372,54404,58042,60874,63187,65140,0),
        (41639,49373,54405,58043,60875,63188,65141,0),
        (41641,49375,54406,58044,60875,63188,65141,0),
        (41644,49376,54407,58044,60876,63189,65142,0),
        (41646,49378,54408,58045,60877,63189,65142,0),
        (41648,49379,54409,58046,60877,63190,65143,0),
        (41651,49381,54410,58047,60878,63190,65143,0),
        (41653,49382,54411,58047,60878,63191,65144,0),
        (41655,49384,54412,58049,60879,63191,65144,0),
        (41657,49386,54413,58049,60880,63192,65144,0),
        (41661,49387,54414,58050,60880,63192,65145,0),
        (41663,49388,54415,58051,60881,63193,65145,0),
        (41665,49389,54416,58052,60882,63193,65146,0),
        (41668,49391,54417,58052,60882,63194,65146,0),
        (41670,49393,54418,58053,60883,63194,65147,0),
        (41672,49394,54419,58054,60883,63195,65147,0),
        (41674,49396,54420,58055,60884,63195,65147,0),
        (41677,49397,54421,58055,60884,63196,65148,0),
        (41679,49399,54422,58056,60885,63197,65148,0),
        (41681,49400,54424,58057,60886,63197,65149,0),
        (41685,49402,54424,58058,60886,63197,65149,0),
        (41687,49403,54425,58058,60887,63198,65150,0),
        (41689,49404,54426,58059,60888,63199,65150,0),
        (41691,49406,54428,58060,60888,63199,65150,0),
        (41694,49408,54428,58061,60889,63199,65151,0),
        (41696,49409,54429,58061,60890,63200,65151,0),
        (41698,49410,54431,58062,60890,63201,65152,0),
        (41701,49412,54432,58063,60891,63201,65152,0),
        (41703,49413,54433,58064,60891,63202,65153,0),
        (41705,49415,54433,58065,60892,63202,65153,0),
        (41707,49417,54435,58065,60893,63203,65154,0),
        (41711,49418,54436,58066,60893,63203,65154,0),
        (41713,49419,54437,58067,60894,63204,65155,0),
        (41715,49421,54438,58068,60895,63204,65155,0),
        (41718,49422,54439,58068,60895,63205,65155,0),
        (41720,49424,54440,58069,60896,63205,65156,0),
        (41722,49425,54441,58070,60896,63206,65156,0),
        (41724,49427,54442,58071,60897,63206,65157,0),
        (41727,49428,54443,58072,60897,63207,65157,0),
        (41729,49430,54444,58072,60898,63207,65158,0),
        (41731,49431,54445,58073,60899,63208,65158,0),
        (41734,49433,54446,58074,60899,63208,65158,0),
        (41737,49434,54447,58075,60900,63209,65159,0),
        (41739,49435,54448,58076,60901,63209,65159,0),
        (41741,49437,54449,58076,60901,63210,65160,0),
        (41744,49439,54450,58077,60902,63210,65160,0),
        (41746,49440,54451,58078,60903,63211,65161,0),
        (41748,49441,54452,58079,60903,63211,65161,0),
        (41751,49443,54453,58079,60904,63212,65161,0),
        (41753,49444,54454,58080,60904,63213,65162,0),
        (41755,49446,54455,58081,60905,63213,65162,0),
        (41757,49448,54456,58082,60906,63213,65163,0),
        (41760,49449,54457,58082,60906,63214,65163,0),
        (41763,49450,54458,58083,60907,63215,65164,0),
        (41765,49452,54459,58084,60908,63215,65164,0),
        (41768,49453,54460,58085,60908,63215,65165,0),
        (41770,49455,54461,58085,60909,63216,65165,0),
        (41772,49456,54462,58086,60909,63217,65166,0),
        (41774,49458,54463,58087,60910,63217,65166,0),
        (41777,49459,54464,58088,60910,63217,65166,0),
        (41779,49461,54465,58088,60911,63218,65167,0),
        (41781,49462,54466,58089,60912,63219,65167,0),
        (41784,49464,54467,58090,60912,63219,65168,0),
        (41786,49465,54468,58091,60913,63220,65168,0),
        (41788,49466,54469,58092,60914,63220,65169,0),
        (41791,49468,54470,58092,60914,63221,65169,0),
        (41794,49470,54471,58093,60915,63221,65170,0),
        (41796,49471,54472,58094,60916,63222,65170,0),
        (41798,49472,54474,58095,60916,63222,65170,0),
        (41801,49474,54474,58095,60917,63223,65171,0),
        (41803,49475,54475,58096,60917,63223,65171,0),
        (41805,49477,54476,58097,60918,63224,65172,0),
        (41807,49479,54478,58098,60919,63224,65172,0),
        (41810,49480,54479,58099,60919,63225,65173,0),
        (41812,49481,54479,58099,60920,63225,65173,0),
        (41814,49482,54481,58100,60920,63226,65173,0),
        (41817,49484,54482,58101,60921,63226,65174,0),
        (41820,49486,54483,58102,60922,63227,65174,0),
        (41822,49487,54483,58103,60922,63227,65175,0),
        (41824,49489,54485,58103,60923,63228,65175,0),
        (41827,49490,54486,58104,60923,63228,65176,0),
        (41829,49491,54487,58105,60924,63229,65176,0),
        (41831,49493,54488,58106,60925,63229,65176,0),
        (41834,49495,54489,58106,60925,63230,65177,0),
        (41836,49496,54490,58107,60926,63231,65177,0),
        (41838,49497,54491,58108,60927,63231,65178,0),
        (41840,49499,54492,58109,60927,63231,65178,0),
        (41843,49500,54493,58109,60928,63232,65179,0),
        (41845,49502,54494,58110,60929,63233,65179,0),
        (41847,49504,54495,58111,60929,63233,65180,0),
        (41851,49505,54496,58112,60930,63233,65180,0),
        (41853,49506,54497,58112,60930,63234,65181,0),
        (41855,49508,54498,58113,60931,63235,65181,0),
        (41858,49509,54499,58114,60932,63235,65181,0),
        (41860,49511,54500,58115,60932,63236,65182,0),
        (41862,49512,54501,58116,60933,63236,65182,0),
        (41864,49514,54502,58116,60933,63237,65183,0),
        (41867,49515,54503,58117,60934,63237,65183,0),
        (41869,49517,54504,58118,60935,63238,65184,0),
        (41871,49518,54505,58119,60935,63238,65184,0),
        (41874,49520,54506,58119,60936,63239,65184,0),
        (41876,49521,54507,58120,60936,63239,65185,0),
        (41878,49522,54508,58121,60937,63240,65185,0),
        (41880,49524,54509,58122,60938,63240,65186,0),
        (41884,49526,54510,58122,60938,63241,65186,0),
        (41886,49527,54511,58123,60939,63241,65187,0),
        (41888,49528,54512,58124,60940,63242,65187,0),
        (41891,49530,54513,58125,60940,63242,65187,0),
        (41893,49531,54514,58125,60941,63243,65188,0),
        (41895,49533,54515,58126,60942,63243,65188,0),
        (41897,49535,54516,58127,60942,63244,65189,0),
        (41900,49536,54517,58128,60943,63244,65189,0),
        (41902,49537,54518,58128,60943,63245,65190,0),
        (41904,49538,54519,58129,60944,63245,65190,0),
        (41907,49540,54520,58130,60945,63246,65191,0),
        (41909,49542,54521,58131,60945,63246,65191,0),
        (41911,49543,54522,58132,60946,63247,65192,0),
        (41913,49545,54523,58133,60946,63247,65192,0),
        (41917,49546,54524,58133,60947,63248,65192,0),
        (41919,49547,54525,58134,60948,63249,65193,0),
        (41921,49549,54527,58135,60948,63249,65193,0),
        (41924,49551,54527,58136,60949,63249,65194,0),
        (41926,49552,54528,58136,60949,63250,65194,0),
        (41928,49553,54529,58137,60950,63251,65195,0),
        (41930,49555,54531,58138,60951,63251,65195,0),
        (41933,49556,54531,58139,60951,63251,65196,0),
        (41935,49558,54532,58139,60952,63252,65196,0),
        (41937,49559,54534,58140,60953,63253,65196,0),
        (41940,49561,54535,58141,60953,63253,65197,0),
        (41942,49562,54535,58142,60954,63254,65197,0),
        (41944,49563,54536,58143,60954,63254,65198,0),
        (41946,49565,54538,58143,60955,63255,65198,0),
        (41950,49567,54539,58144,60956,63255,65199,0),
        (41952,49568,54539,58145,60956,63256,65199,0),
        (41954,49569,54541,58146,60957,63256,65199,0),
        (41957,49571,54542,58146,60957,63257,65200,0),
        (41959,49572,54543,58147,60958,63257,65200,0),
        (41961,49574,54543,58148,60959,63258,65201,0),
        (41963,49576,54545,58149,60959,63258,65201,0),
        (41966,49577,54546,58149,60960,63259,65202,0),
        (41968,49578,54547,58150,60961,63259,65202,0),
        (41970,49579,54548,58151,60961,63260,65202,0),
        (41973,49581,54549,58152,60962,63260,65203,0),
        (41975,49583,54550,58152,60962,63261,65203,0),
        (41977,49584,54551,58153,60963,63261,65204,0),
        (41979,49586,54552,58154,60964,63262,65204,0),
        (41982,49587,54553,58155,60964,63262,65205,0),
        (41984,49588,54554,58155,60965,63263,65205,0),
        (41986,49590,54555,58156,60966,63263,65206,0),
        (41990,49591,54556,58157,60966,63264,65206,0),
        (41992,49593,54557,58158,60967,63264,65207,0),
        (41994,49594,54558,58159,60967,63265,65207,0),
        (41996,49596,54559,58159,60968,63265,65207,0),
        (41999,49597,54560,58160,60968,63266,65208,0),
        (42001,49599,54561,58161,60969,63266,65208,0),
        (42003,49600,54562,58162,60970,63267,65209,0),
        (42006,49602,54563,58162,60970,63267,65209,0),
        (42008,49603,54564,58163,60971,63268,65210,0),
        (42010,49604,54565,58164,60972,63268,65210,0),
        (42012,49606,54566,58165,60972,63269,65210,0),
        (42015,49607,54567,58165,60973,63269,65211,0),
        (42017,49609,54568,58166,60974,63270,65211,0),
        (42019,49610,54569,58167,60974,63271,65212,0),
        (42022,49612,54570,58168,60975,63271,65212,0),
        (42024,49613,54571,58168,60975,63272,65213,0),
        (42026,49614,54572,58169,60976,63272,65213,0),
        (42029,49616,54573,58170,60977,63273,65213,0),
        (42032,49618,54574,58171,60977,63273,65214,0),
        (42034,49619,54575,58171,60978,63274,65214,0),
        (42036,49620,54576,58172,60978,63274,65215,0),
        (42039,49622,54577,58173,60979,63275,65215,0),
        (42041,49623,54578,58174,60980,63275,65216,0),
        (42043,49625,54579,58175,60980,63276,65216,0),
        (42045,49627,54580,58175,60981,63276,65216,0),
        (42048,49628,54581,58176,60981,63277,65217,0),
        (42050,49629,54582,58177,60982,63277,65217,0),
        (42052,49630,54583,58178,60983,63278,65218,0),
        (42055,49632,54584,58179,60983,63278,65218,0),
        (42057,49634,54585,58179,60984,63279,65219,0),
        (42059,49635,54586,58180,60985,63279,65219,0),
        (42061,49637,54587,58181,60985,63280,65220,0),
        (42064,49638,54588,58182,60986,63280,65220,0),
        (42066,49639,54589,58182,60986,63281,65221,0),
        (42068,49641,54590,58183,60987,63281,65221,0),
        (42072,49642,54591,58184,60988,63282,65221,0),
        (42074,49644,54592,58185,60988,63282,65222,0),
        (42076,49645,54593,58186,60989,63283,65222,0),
        (42078,49647,54594,58186,60989,63283,65223,0),
        (42081,49648,54595,58187,60990,63284,65223,0),
        (42083,49649,54596,58188,60991,63284,65224,0),
        (42085,49651,54597,58189,60991,63285,65224,0),
        (42088,49653,54598,58189,60992,63285,65224,0),
        (42090,49654,54599,58190,60992,63286,65225,0),
        (42092,49655,54600,58191,60993,63286,65225,0),
        (42094,49657,54601,58192,60994,63287,65226,0),
        (42097,49658,54602,58192,60994,63287,65226,0),
        (42099,49660,54603,58193,60995,63288,65227,0),
        (42101,49661,54604,58194,60996,63288,65227,0),
        (42104,49663,54605,58195,60996,63289,65227,0),
        (42106,49664,54606,58195,60997,63290,65228,0),
        (42108,49665,54607,58196,60998,63290,65228,0),
        (42110,49667,54608,58197,60998,63290,65229,0),
        (42113,49669,54609,58198,60999,63291,65229,0),
        (42115,49670,54610,58198,60999,63292,65230,0),
        (42117,49671,54612,58199,61000,63292,65230,0),
        (42120,49673,54612,58200,61000,63292,65230,0),
        (42123,49674,54613,58201,61001,63293,65231,0),
        (42125,49676,54614,58202,61002,63294,65231,0),
        (42127,49677,54616,58202,61002,63294,65232,0),
        (42130,49679,54616,58203,61003,63294,65232,0),
        (42132,49680,54617,58204,61004,63295,65233,0),
        (42134,49681,54619,58205,61004,63296,65233,0),
        (42137,49683,54619,58205,61005,63296,65234,0),
        (42139,49684,54620,58206,61005,63297,65234,0),
        (42141,49686,54621,58207,61006,63297,65235,0),
        (42143,49688,54623,58208,61007,63298,65235,0),
        (42146,49689,54623,58208,61007,63298,65235,0),
        (42148,49690,54624,58209,61008,63299,65236,0),
        (42150,49691,54626,58210,61009,63299,65236,0),
        (42153,49693,54627,58211,61009,63300,65237,0),
        (42155,49695,54627,58211,61010,63300,65237,0),
        (42157,49696,54628,58212,61010,63301,65238,0),
        (42159,49698,54630,58213,61011,63301,65238,0),
        (42162,49699,54631,58214,61011,63302,65239,0),
        (42164,49700,54631,58214,61012,63302,65239,0),
        (42166,49702,54633,58215,61013,63303,65239,0),
        (42169,49703,54634,58216,61013,63303,65240,0),
        (42171,49705,54634,58217,61014,63304,65240,0),
        (42173,49706,54635,58218,61015,63304,65241,0),
        (42175,49708,54637,58218,61015,63305,65241,0),
        (42179,49709,54638,58219,61016,63305,65242,0),
        (42181,49710,54638,58220,61017,63306,65242,0),
        (42183,49712,54640,58221,61017,63306,65242,0),
        (42186,49714,54641,58221,61018,63307,65243,0),
        (42188,49715,54642,58222,61018,63307,65243,0),
        (42190,49716,54642,58223,61019,63308,65244,0),
        (42192,49718,54644,58224,61020,63308,65244,0),
        (42195,49719,54645,58224,61020,63309,65245,0),
        (42197,49721,54645,58225,61021,63309,65245,0),
        (42199,49722,54647,58226,61021,63310,65245,0),
        (42202,49724,54648,58227,61022,63310,65246,0),
        (42204,49725,54649,58227,61022,63311,65246,0),
        (42206,49726,54649,58228,61023,63311,65247,0),
        (42208,49728,54651,58229,61024,63312,65247,0),
        (42211,49729,54652,58230,61024,63312,65248,0),
        (42213,49731,54653,58230,61025,63313,65248,0),
        (42215,49732,54654,58231,61026,63313,65249,0),
        (42218,49734,54655,58232,61026,63314,65249,0),
        (42220,49735,54656,58233,61027,63315,65249,0),
        (42222,49736,54656,58234,61028,63315,65250,0),
        (42224,49738,54658,58234,61028,63316,65250,0),
        (42227,49740,54659,58235,61029,63316,65251,0),
        (42229,49741,54660,58236,61029,63317,65251,0),
        (42231,49742,54661,58237,61030,63317,65252,0),
        (42234,49744,54662,58237,61030,63318,65252,0),
        (42236,49745,54663,58238,61031,63318,65253,0),
        (42238,49747,54664,58239,61032,63319,65253,0),
        (42240,49748,54665,58240,61032,63319,65253,0),
        (42243,49750,54666,58240,61033,63320,65254,0),
        (42245,49751,54667,58241,61034,63320,65254,0),
        (42247,49752,54668,58242,61034,63321,65255,0),
        (42251,49754,54669,58243,61035,63321,65255,0),
        (42253,49755,54670,58243,61035,63322,65256,0),
        (42255,49757,54671,58244,61036,63322,65256,0),
        (42257,49759,54672,58245,61037,63323,65256,0),
        (42260,49760,54673,58246,61037,63323,65257,0),
        (42262,49761,54674,58246,61038,63324,65257,0),
        (42264,49762,54675,58247,61039,63324,65258,0),
        (42267,49764,54676,58248,61039,63325,65258,0),
        (42269,49765,54677,58249,61040,63325,65259,0),
        (42271,49767,54678,58250,61040,63326,65259,0),
        (42273,49769,54679,58250,61041,63326,65259,0),
        (42276,49770,54680,58251,61041,63327,65260,0),
        (42278,49771,54681,58252,61042,63327,65260,0),
        (42280,49772,54682,58253,61043,63328,65261,0),
        (42283,49774,54683,58253,61043,63328,65261,0),
        (42285,49776,54684,58254,61044,63329,65262,0),
        (42287,49777,54685,58255,61045,63329,65262,0),
        (42289,49779,54686,58256,61045,63330,65262,0),
        (42292,49780,54687,58256,61046,63330,65263,0),
        (42294,49781,54688,58257,61047,63331,65263,0),
        (42296,49782,54689,58258,61047,63331,65264,0),
        (42299,49784,54690,58259,61048,63332,65264,0),
        (42301,49786,54691,58259,61048,63332,65265,0),
        (42303,49787,54692,58260,61049,63333,65265,0),
        (42305,49789,54693,58261,61049,63333,65266,0),
        (42308,49790,54694,58262,61050,63334,65266,0),
        (42310,49791,54695,58262,61051,63334,65267,0),
        (42312,49793,54696,58263,61051,63335,65267,0),
        (42315,49794,54697,58264,61052,63335,65267,0),
        (42317,49796,54698,58265,61052,63336,65268,0),
        (42319,49797,54699,58266,61053,63336,65268,0),
        (42321,49799,54700,58266,61054,63337,65269,0),
        (42324,49800,54701,58267,61054,63337,65269,0),
        (42326,49801,54702,58268,61055,63338,65270,0),
        (42328,49803,54703,58269,61056,63338,65270,0),
        (42331,49805,54704,58269,61056,63339,65270,0),
        (42333,49806,54705,58270,61057,63340,65271,0),
        (42335,49807,54706,58271,61058,63340,65271,0),
        (42337,49809,54707,58272,61058,63341,65272,0),
        (42340,49810,54708,58272,61059,63341,65272,0),
        (42342,49811,54709,58273,61059,63342,65273,0),
        (42344,49813,54710,58274,61060,63342,65273,0),
        (42347,49815,54711,58275,61060,63343,65273,0),
        (42349,49816,54712,58275,61061,63343,65274,0),
        (42352,49817,54713,58276,61062,63344,65274,0),
        (42354,49819,54714,58277,61062,63344,65275,0),
        (42357,49820,54715,58278,61063,63345,65275,0),
        (42359,49821,54716,58278,61064,63345,65276,0),
        (42361,49823,54717,58279,61064,63346,65276,0),
        (42364,49825,54718,58280,61065,63346,65276,0),
        (42366,49826,54719,58281,61065,63347,65277,0),
        (42368,49827,54720,58282,61066,63347,65277,0),
        (42370,49829,54721,58282,61067,63348,65278,0),
        (42373,49830,54722,58283,61067,63348,65278,0),
        (42375,49832,54723,58284,61068,63349,65279,0),
        (42377,49833,54724,58285,61068,63349,65279,0),
        (42380,49835,54725,58285,61069,63350,65280,0),
        (42382,49836,54726,58286,61070,63350,65280,0),
        (42384,49837,54727,58287,61070,63351,65280,0),
        (42386,49839,54728,58288,61071,63351,65281,0),
        (42389,49840,54729,58288,61071,63352,65281,0),
        (42391,49842,54730,58289,61072,63352,65282,0),
        (42393,49843,54731,58290,61073,63353,65282,0),
        (42396,49845,54732,58291,61073,63353,65283,0),
        (42398,49846,54733,58291,61074,63354,65283,0),
        (42400,49847,54734,58292,61075,63354,65284,0),
        (42402,49849,54735,58293,61075,63355,65284,0),
        (42405,49850,54736,58294,61076,63355,65284,0),
        (42407,49852,54737,58294,61076,63356,65285,0),
        (42409,49853,54738,58295,61077,63356,65285,0),
        (42412,49855,54739,58296,61078,63357,65286,0),
        (42414,49856,54740,58297,61078,63357,65286,0),
        (42416,49857,54741,58298,61079,63358,65287,0),
        (42418,49859,54742,58298,61079,63358,65287,0),
        (42421,49860,54743,58299,61080,63359,65288,0),
        (42423,49862,54744,58300,61081,63359,65288,0),
        (42425,49863,54745,58301,61081,63360,65288,0),
        (42428,49865,54746,58301,61082,63360,65289,0),
        (42430,49866,54747,58302,61082,63361,65289,0),
        (42432,49867,54748,58303,61083,63361,65290,0),
        (42434,49869,54749,58304,61084,63362,65290,0),
        (42437,49870,54750,58304,61084,63362,65291,0),
        (42439,49872,54751,58305,61085,63363,65291,0),
        (42441,49873,54752,58306,61086,63363,65291,0),
        (42444,49875,54753,58307,61086,63364,65292,0),
        (42446,49876,54754,58307,61087,63365,65292,0),
        (42448,49877,54755,58308,61087,63365,65293,0),
        (42450,49879,54756,58309,61088,63365,65293,0),
        (42453,49880,54757,58310,61088,63366,65294,0),
        (42455,49882,54758,58310,61089,63367,65294,0),
        (42457,49883,54759,58311,61090,63367,65294,0),
        (42460,49885,54760,58312,61090,63367,65295,0),
        (42462,49886,54761,58313,61091,63368,65295,0),
        (42464,49887,54762,58314,61092,63369,65296,0),
        (42466,49889,54763,58314,61092,63369,65296,0),
        (42469,49890,54764,58315,61093,63369,65297,0),
        (42471,49892,54765,58316,61094,63370,65297,0),
        (42473,49893,54766,58316,61094,63371,65297,0),
        (42476,49895,54767,58317,61095,63371,65298,0),
        (42478,49896,54768,58318,61095,63372,65298,0),
        (42480,49897,54769,58319,61096,63372,65299,0),
        (42483,49899,54770,58319,61096,63373,65299,0),
        (42485,49900,54771,58320,61097,63373,65300,0),
        (42487,49902,54772,58321,61098,63374,65300,0),
        (42489,49904,54773,58322,61098,63374,65301,0),
        (42492,49905,54774,58322,61099,63375,65301,0),
        (42494,49906,54775,58323,61100,63375,65301,0),
        (42496,49907,54776,58324,61100,63376,65302,0),
        (42499,49909,54777,58325,61101,63376,65302,0),
        (42501,49910,54778,58325,61101,63377,65303,0),
        (42503,49912,54779,58326,61102,63377,65303,0),
        (42505,49914,54780,58327,61103,63378,65304,0),
        (42508,49915,54781,58328,61103,63378,65304,0),
        (42510,49916,54782,58328,61104,63379,65305,0),
        (42512,49917,54783,58329,61104,63379,65305,0),
        (42515,49919,54784,58330,61105,63380,65305,0),
        (42517,49920,54785,58331,61106,63380,65306,0),
        (42519,49922,54786,58332,61106,63381,65306,0),
        (42521,49924,54787,58332,61107,63381,65307,0),
        (42524,49925,54788,58333,61107,63382,65307,0),
        (42526,49926,54789,58334,61108,63382,65308,0),
        (42528,49927,54790,58335,61109,63383,65308,0),
        (42531,49929,54791,58335,61109,63383,65308,0),
        (42533,49930,54792,58336,61110,63384,65309,0),
        (42535,49932,54793,58337,61111,63384,65309,0),
        (42537,49934,54794,58338,61111,63385,65310,0),
        (42540,49935,54795,58338,61112,63385,65310,0),
        (42542,49936,54796,58339,61112,63386,65311,0),
        (42544,49937,54797,58340,61113,63386,65311,0),
        (42547,49939,54798,58341,61114,63387,65311,0),
        (42549,49940,54799,58341,61114,63387,65312,0),
        (42551,49942,54800,58342,61115,63388,65312,0),
        (42553,49944,54801,58343,61115,63388,65313,0),
        (42556,49945,54802,58344,61116,63389,65313,0),
        (42558,49946,54803,58344,61117,63389,65314,0),
        (42560,49947,54804,58345,61117,63390,65314,0),
        (42563,49949,54805,58346,61118,63390,65314,0),
        (42565,49950,54806,58347,61118,63391,65315,0),
        (42567,49952,54806,58348,61119,63391,65315,0),
        (42569,49953,54808,58348,61120,63392,65316,0),
        (42572,49955,54809,58349,61120,63392,65316,0),
        (42574,49956,54810,58350,61121,63393,65317,0),
        (42576,49957,54811,58351,61121,63393,65317,0),
        (42579,49959,54812,58351,61122,63394,65317,0),
        (42581,49960,54813,58352,61123,63395,65318,0),
        (42583,49962,54813,58353,61123,63395,65318,0),
        (42585,49963,54815,58354,61124,63395,65319,0),
        (42588,49965,54816,58354,61124,63396,65319,0),
        (42590,49966,54816,58355,61125,63397,65320,0),
        (42592,49967,54818,58356,61126,63397,65320,0),
        (42595,49969,54819,58357,61126,63397,65321,0),
        (42597,49970,54820,58357,61127,63398,65321,0),
        (42599,49972,54820,58358,61128,63399,65321,0),
        (42601,49973,54822,58359,61128,63399,65322,0),
        (42604,49975,54823,58360,61129,63399,65322,0),
        (42606,49976,54823,58360,61129,63400,65323,0),
        (42608,49977,54825,58361,61130,63401,65323,0),
        (42611,49979,54826,58362,61131,63401,65324,0),
        (42613,49980,54826,58362,61131,63402,65324,0),
        (42615,49981,54827,58363,61132,63402,65325,0),
        (42617,49983,54829,58364,61132,63403,65325,0),
        (42620,49985,54829,58365,61133,63403,65325,0),
        (42622,49986,54830,58365,61134,63404,65326,0),
        (42624,49987,54832,58366,61134,63404,65326,0),
        (42626,49989,54833,58367,61135,63405,65327,0),
        (42628,49990,54833,58368,61135,63405,65327,0),
        (42630,49991,54834,58369,61136,63406,65328,0),
        (42632,49993,54836,58369,61137,63406,65328,0),
        (42635,49995,54836,58370,61137,63407,65329,0),
        (42637,49996,54837,58371,61138,63407,65329,0),
        (42639,49997,54839,58372,61138,63408,65329,0),
        (42642,49999,54839,58372,61139,63408,65330,0),
        (42644,50000,54840,58373,61140,63409,65330,0),
        (42646,50001,54841,58374,61140,63409,65331,0),
        (42648,50003,54843,58375,61141,63410,65331,0),
        (42651,50004,54843,58375,61141,63410,65332,0),
        (42653,50006,54844,58376,61142,63411,65332,0),
        (42655,50007,54846,58377,61143,63411,65332,0),
        (42658,50009,54846,58378,61143,63412,65333,0),
        (42660,50010,54847,58378,61144,63412,65333,0),
        (42662,50011,54848,58379,61145,63413,65334,0),
        (42664,50013,54849,58380,61145,63413,65334,0),
        (42667,50014,54850,58381,61146,63414,65335,0),
        (42669,50016,54851,58381,61146,63414,65335,0),
        (42671,50017,54852,58382,61147,63415,65335,0),
        (42674,50019,54853,58383,61148,63415,65336,0),
        (42676,50020,54854,58384,61148,63416,65336,0),
        (42678,50021,54855,58385,61149,63416,65337,0),
        (42680,50023,54856,58385,61149,63417,65337,0),
        (42683,50024,54857,58386,61150,63417,65338,0),
        (42685,50026,54858,58387,61151,63418,65338,0),
        (42687,50027,54859,58388,61151,63418,65338,0),
        (42690,50029,54860,58388,61152,63419,65339,0),
        (42692,50030,54861,58389,61152,63419,65339,0),
        (42694,50031,54862,58390,61153,63420,65340,0),
        (42696,50033,54863,58391,61154,63420,65340,0),
        (42699,50034,54864,58391,61154,63421,65341,0),
        (42701,50035,54865,58392,61155,63421,65341,0),
        (42703,50037,54866,58393,61155,63422,65341,0),
        (42706,50039,54867,58394,61156,63422,65342,0),
        (42708,50040,54868,58394,61157,63423,65342,0),
        (42710,50041,54869,58395,61157,63423,65343,0),
        (42712,50043,54870,58396,61158,63424,65343,0),
        (42715,50044,54871,58396,61158,63424,65344,0),
        (42717,50045,54872,58397,61159,63425,65344,0),
        (42719,50047,54873,58398,61160,63425,65344,0),
        (42722,50048,54874,58399,61160,63426,65345,0),
        (42724,50050,54875,58399,61161,63427,65345,0),
        (42725,50051,54876,58400,61162,63427,65346,0),
        (42727,50053,54877,58401,61162,63427,65346,0),
        (42730,50054,54878,58402,61163,63428,65347,0),
        (42732,50055,54879,58402,61163,63428,65347,0),
        (42734,50056,54880,58403,61164,63429,65348,0),
        (42737,50058,54881,58404,61164,63429,65348,0),
        (42739,50060,54882,58405,61165,63430,65348,0),
        (42741,50061,54883,58406,61166,63430,65349,0),
        (42743,50063,54884,58406,61166,63431,65349,0),
        (42746,50064,54885,58407,61167,63431,65350,0),
        (42748,50065,54886,58408,61168,63432,65350,0),
        (42750,50066,54887,58409,61168,63432,65351,0),
        (42753,50068,54888,58409,61169,63433,65351,0),
        (42755,50069,54889,58410,61169,63434,65352,0),
        (42757,50071,54890,58411,61170,63434,65352,0),
        (42759,50073,54891,58412,61171,63434,65352,0),
        (42762,50074,54892,58412,61171,63435,65353,0),
        (42764,50075,54893,58413,61172,63436,65353,0),
        (42766,50076,54894,58414,61172,63436,65354,0),
        (42769,50078,54895,58415,61173,63436,65354,0),
        (42771,50079,54896,58415,61173,63437,65355,0),
        (42773,50081,54897,58416,61174,63438,65355,0),
        (42775,50082,54898,58417,61175,63438,65355,0),
        (42778,50084,54899,58418,61175,63438,65356,0),
        (42780,50085,54900,58418,61176,63439,65356,0),
        (42782,50086,54901,58419,61177,63440,65357,0),
        (42785,50088,54902,58420,61177,63440,65357,0),
        (42787,50089,54903,58420,61178,63441,65358,0),
        (42789,50090,54903,58421,61179,63441,65358,0),
        (42791,50092,54905,58422,61179,63442,65358,0),
        (42793,50094,54906,58423,61180,63442,65359,0),
        (42795,50095,54907,58423,61180,63443,65359,0),
        (42797,50096,54908,58424,61181,63443,65360,0),
        (42800,50098,54909,58425,61181,63444,65360,0),
        (42802,50099,54910,58426,61182,63444,65361,0),
        (42804,50100,54910,58427,61183,63445,65361,0),
        (42806,50102,54912,58427,61183,63445,65361,0),
        (42809,50103,54913,58428,61184,63446,65362,0),
        (42811,50105,54913,58429,61185,63446,65362,0),
        (42813,50106,54915,58430,61185,63447,65363,0),
        (42816,50108,54916,58430,61186,63447,65363,0),
        (42818,50109,54916,58431,61186,63448,65364,0),
        (42820,50110,54917,58432,61187,63448,65364,0),
        (42822,50112,54919,58433,61188,63449,65364,0),
        (42825,50113,54919,58433,61188,63449,65365,0),
        (42827,50114,54920,58434,61189,63450,65365,0),
        (42829,50116,54922,58435,61189,63450,65366,0),
        (42832,50118,54922,58436,61190,63451,65366,0),
        (42834,50119,54923,58436,61190,63451,65367,0),
        (42836,50120,54924,58437,61191,63452,65367,0),
        (42838,50122,54925,58438,61192,63452,65367,0),
        (42841,50123,54926,58439,61192,63453,65368,0),
        (42843,50124,54927,58439,61193,63453,65368,0),
        (42845,50126,54928,58440,61194,63454,65369,0),
        (42848,50127,54929,58441,61194,63454,65369,0),
        (42849,50129,54930,58442,61195,63455,65370,0),
        (42851,50130,54931,58443,61195,63455,65370,0),
        (42853,50132,54932,58443,61196,63456,65370,0),
        (42856,50133,54933,58444,61197,63456,65371,0),
        (42858,50134,54934,58444,61197,63457,65371,0),
        (42860,50135,54935,58445,61198,63457,65372,0),
        (42863,50137,54936,58446,61198,63458,65372,0),
        (42865,50138,54937,58447,61199,63458,65373,0),
        (42867,50140,54938,58448,61200,63459,65373,0),
        (42869,50142,54939,58448,61200,63459,65374,0),
        (42872,50143,54940,58449,61201,63460,65374,0),
        (42874,50144,54941,58450,61202,63460,65374,0),
        (42876,50145,54942,58451,61202,63461,65375,0),
        (42879,50147,54943,58451,61203,63461,65375,0),
        (42881,50148,54944,58452,61203,63462,65376,0),
        (42883,50149,54945,58453,61204,63462,65376,0),
        (42885,50151,54946,58454,61204,63463,65377,0),
        (42888,50153,54947,58454,61205,63463,65377,0),
        (42890,50154,54948,58455,61206,63464,65378,0),
        (42892,50155,54949,58456,61206,63464,65378,0),
        (42895,50157,54950,58457,61207,63465,65378,0),
        (42897,50158,54951,58457,61207,63465,65379,0),
        (42898,50159,54952,58458,61208,63466,65379,0),
        (42900,50161,54953,58459,61209,63466,65380,0),
        (42903,50162,54954,58460,61209,63467,65380,0),
        (42905,50164,54955,58460,61210,63467,65381,0),
        (42907,50165,54956,58461,61211,63468,65381,0),
        (42910,50167,54957,58462,61211,63468,65381,0),
        (42912,50168,54958,58463,61212,63469,65382,0),
        (42914,50169,54959,58463,61212,63469,65382,0),
        (42916,50171,54960,58464,61213,63470,65383,0),
        (42919,50172,54961,58465,61213,63470,65383,0),
        (42921,50173,54962,58465,61214,63471,65384,0),
        (42923,50175,54963,58466,61215,63471,65384,0),
        (42926,50176,54964,58467,61215,63472,65384,0),
        (42928,50178,54965,58468,61216,63472,65385,0),
        (42930,50179,54965,58469,61217,63473,65385,0),
        (42932,50181,54967,58469,61217,63473,65386,0),
        (42935,50182,54968,58470,61218,63474,65386,0),
        (42937,50183,54968,58471,61218,63474,65387,0),
        (42939,50184,54970,58472,61219,63475,65387,0),
        (42941,50186,54971,58472,61219,63475,65387,0),
        (42943,50188,54972,58473,61220,63476,65388,0),
        (42945,50189,54972,58474,61221,63476,65388,0),
        (42947,50191,54974,58475,61221,63477,65389,0),
        (42950,50192,54975,58475,61222,63477,65389,0),
        (42952,50193,54975,58476,61223,63478,65390,0),
        (42954,50194,54977,58477,61223,63478,65390,0),
        (42957,50196,54978,58478,61224,63479,65390,0),
        (42959,50197,54978,58478,61224,63480,65391,0),
        (42961,50199,54979,58479,61225,63480,65391,0),
        (42963,50200,54981,58480,61226,63480,65392,0),
        (42966,50202,54981,58481,61226,63481,65392,0),
        (42968,50203,54982,58481,61227,63482,65393,0),
        (42970,50204,54984,58482,61227,63482,65393,0),
        (42973,50206,54984,58483,61228,63482,65393,0),
        (42975,50207,54985,58483,61228,63483,65394,0),
        (42977,50208,54986,58484,61229,63484,65394,0),
        (42978,50210,54987,58485,61230,63484,65395,0),
        (42981,50211,54988,58486,61230,63484,65395,0),
        (42983,50213,54989,58486,61231,63485,65396,0),
        (42985,50214,54990,58487,61232,63485,65396,0),
        (42988,50216,54991,58488,61232,63486,65396,0),
        (42990,50217,54992,58489,61233,63487,65397,0),
        (42992,50218,54993,58490,61233,63487,65397,0),
        (42994,50220,54994,58490,61234,63487,65398,0),
        (42997,50221,54995,58491,61235,63488,65398,0),
        (42999,50222,54996,58492,61235,63489,65399,0),
        (43001,50224,54997,58493,61236,63489,65399,0),
        (43004,50225,54998,58493,61236,63489,65399,0),
        (43006,50227,54999,58494,61237,63490,65400,0),
        (43008,50228,55000,58495,61238,63491,65400,0),
        (43010,50230,55001,58496,61238,63491,65401,0),
        (43013,50231,55002,58496,61239,63491,65401,0),
        (43014,50232,55003,58497,61240,63492,65402,0),
        (43016,50233,55004,58498,61240,63493,65402,0),
        (43019,50235,55005,58499,61241,63493,65403,0),
        (43021,50236,55006,58499,61241,63494,65403,0),
        (43023,50238,55007,58500,61242,63494,65403,0),
        (43025,50239,55008,58501,61242,63495,65404,0),
        (43028,50241,55009,58501,61243,63495,65404,0),
        (43030,50242,55010,58502,61244,63496,65405,0),
        (43032,50243,55011,58503,61244,63496,65405,0),
        (43035,50245,55012,58504,61245,63497,65406,0),
        (43037,50246,55013,58504,61245,63497,65406,0),
        (43039,50247,55014,58505,61246,63498,65406,0),
        (43041,50249,55015,58506,61247,63498,65407,0),
        (43044,50250,55016,58507,61247,63498,65407,0),
        (43046,50252,55017,58507,61248,63499,65408,0),
        (43048,50253,55018,58508,61248,63500,65408,0),
        (43050,50255,55019,58509,61249,63500,65409,0),
        (43052,50256,55019,58510,61250,63501,65409,0),
        (43054,50257,55020,58511,61250,63501,65410,0),
        (43056,50259,55022,58511,61251,63502,65410,0),
        (43059,50260,55022,58512,61251,63502,65410,0),
        (43061,50261,55023,58513,61252,63503,65411,0),
        (43063,50263,55025,58514,61253,63503,65411,0),
        (43066,50264,55025,58514,61253,63504,65412,0),
        (43068,50266,55026,58515,61254,63504,65412,0),
        (43070,50267,55027,58516,61255,63505,65413,0),
        (43072,50269,55028,58516,61255,63505,65413,0),
        (43075,50270,55029,58517,61256,63506,65413,0),
        (43077,50271,55030,58518,61256,63506,65414,0),
        (43079,50272,55031,58519,61257,63507,65414,0),
        (43081,50274,55032,58519,61257,63507,65415,0),
        (43083,50275,55033,58520,61258,63508,65415,0),
        (43085,50277,55034,58521,61259,63508,65416,0),
        (43087,50278,55035,58522,61259,63509,65416,0),
        (43090,50280,55036,58522,61260,63509,65417,0),
        (43092,50281,55037,58523,61261,63510,65417,0),
        (43094,50282,55038,58524,61261,63510,65417,0),
        (43097,50284,55039,58525,61262,63511,65418,0),
        (43099,50285,55040,58525,61262,63511,65418,0),
        (43101,50286,55041,58526,61263,63512,65419,0),
        (43104,50288,55042,58527,61263,63512,65419,0),
        (43106,50289,55043,58528,61264,63513,65420,0),
        (43108,50291,55044,58529,61265,63513,65420,0),
        (43110,50292,55045,58529,61265,63514,65420,0),
        (43112,50294,55046,58530,61266,63514,65421,0),
        (43114,50295,55047,58531,61267,63515,65421,0),
        (43116,50296,55048,58531,61267,63515,65422,0),
        (43119,50298,55049,58532,61268,63516,65422,0),
        (43121,50299,55050,58533,61268,63516,65423,0),
        (43123,50300,55051,58534,61269,63517,65423,0),
        (43125,50302,55052,58534,61270,63517,65423,0),
        (43128,50303,55053,58535,61270,63518,65424,0),
        (43130,50305,55054,58536,61271,63518,65424,0),
        (43132,50306,55055,58537,61271,63519,65425,0),
        (43135,50308,55056,58537,61272,63519,65425,0),
        (43137,50309,55057,58538,61272,63520,65426,0),
        (43138,50310,55058,58539,61273,63520,65426,0),
        (43140,50312,55059,58540,61274,63521,65426,0),
        (43143,50313,55060,58540,61274,63521,65427,0),
        (43145,50314,55060,58541,61275,63522,65427,0),
        (43147,50316,55062,58542,61276,63522,65428,0),
        (43150,50317,55063,58543,61276,63523,65428,0),
        (43152,50319,55063,58543,61277,63523,65429,0),
        (43154,50320,55064,58544,61277,63524,65429,0),
        (43156,50322,55066,58545,61278,63524,65429,0),
        (43159,50323,55066,58545,61278,63525,65430,0),
        (43161,50324,55067,58546,61279,63525,65430,0),
        (43163,50325,55069,58547,61280,63526,65431,0),
        (43166,50327,55069,58548,61280,63526,65431,0),
        (43167,50328,55070,58548,61281,63527,65432,0),
        (43169,50329,55071,58549,61282,63527,65432,0),
        (43171,50331,55072,58550,61282,63528,65432,0),
        (43174,50332,55073,58551,61283,63528,65433,0),
        (43176,50334,55074,58551,61283,63529,65433,0),
        (43178,50335,55075,58552,61284,63529,65434,0),
        (43181,50337,55076,58553,61284,63530,65434,0),
        (43183,50338,55077,58554,61285,63530,65435,0),
        (43185,50339,55078,58555,61286,63531,65435,0),
        (43187,50341,55079,58555,61286,63531,65435,0),
        (43190,50342,55080,58556,61287,63532,65436,0),
        (43192,50343,55081,58557,61288,63532,65436,0),
        (43193,50345,55082,58558,61288,63533,65437,0),
        (43196,50346,55083,58558,61289,63533,65437,0),
        (43198,50348,55084,58559,61289,63534,65438,0),
        (43200,50349,55085,58560,61290,63534,65438,0),
        (43202,50351,55086,58560,61291,63535,65438,0),
        (43205,50352,55087,58561,61291,63535,65439,0),
        (43207,50353,55088,58562,61292,63536,65439,0),
        (43209,50354,55089,58563,61292,63536,65440,0),
        (43212,50356,55090,58563,61293,63537,65440,0),
        (43214,50357,55091,58564,61293,63537,65441,0),
        (43216,50359,55092,58565,61294,63538,65441,0),
        (43217,50360,55093,58566,61295,63538,65441,0),
        (43220,50362,55094,58566,61295,63539,65442,0),
        (43222,50363,55095,58567,61296,63539,65442,0),
        (43224,50364,55096,58568,61297,63540,65443,0),
        (43227,50366,55097,58569,61297,63540,65443,0),
        (43229,50367,55098,58569,61298,63541,65444,0),
        (43231,50368,55098,58570,61298,63541,65444,0),
        (43233,50370,55100,58571,61299,63542,65444,0),
        (43236,50371,55101,58572,61299,63542,65445,0),
        (43238,50372,55101,58572,61300,63543,65445,0),
        (43240,50374,55103,58573,61301,63543,65446,0),
        (43242,50375,55103,58574,61301,63544,65446,0),
        (43244,50377,55104,58574,61302,63544,65447,0),
        (43246,50378,55105,58575,61303,63545,65447,0),
        (43248,50380,55106,58576,61303,63545,65447,0),
        (43251,50381,55107,58577,61304,63546,65448,0),
        (43253,50382,55108,58577,61304,63546,65448,0),
        (43255,50383,55109,58578,61305,63547,65449,0),
        (43258,50385,55110,58579,61305,63547,65449,0),
        (43260,50386,55111,58580,61306,63548,65450,0),
        (43262,50388,55112,58581,61307,63548,65450,0),
        (43264,50389,55113,58581,61307,63549,65450,0),
        (43266,50391,55114,58582,61308,63549,65451,0),
        (43268,50392,55115,58583,61309,63550,65451,0),
        (43270,50393,55116,58584,61309,63550,65452,0),
        (43273,50395,55117,58584,61310,63551,65452,0),
        (43275,50396,55118,58585,61310,63551,65453,0),
        (43277,50397,55119,58586,61311,63552,65453,0),
        (43279,50399,55120,58586,61312,63552,65453,0),
        (43282,50400,55121,58587,61312,63553,65454,0),
        (43284,50401,55122,58588,61313,63553,65454,0),
        (43286,50403,55123,58589,61313,63554,65455,0),
        (43288,50404,55124,58589,61314,63554,65455,0),
        (43290,50406,55125,58590,61314,63555,65456,0),
        (43292,50407,55126,58591,61315,63555,65456,0),
        (43294,50409,55127,58592,61316,63556,65457,0),
        (43297,50410,55128,58592,61316,63556,65457,0),
        (43299,50411,55129,58593,61317,63557,65457,0),
        (43301,50412,55130,58594,61318,63557,65458,0),
        (43304,50414,55131,58595,61318,63558,65458,0),
        (43306,50415,55132,58595,61319,63558,65459,0),
        (43308,50416,55132,58596,61319,63559,65459,0),
        (43310,50418,55134,58597,61320,63559,65460,0),
        (43312,50419,55134,58597,61320,63560,65460,0),
        (43314,50421,55135,58598,61321,63560,65460,0),
        (43316,50422,55137,58599,61322,63561,65461,0),
        (43319,50424,55137,58600,61322,63561,65461,0),
        (43321,50425,55138,58600,61323,63562,65462,0),
        (43323,50426,55139,58601,61324,63562,65462,0),
        (43325,50428,55140,58602,61324,63563,65463,0),
        (43328,50429,55141,58603,61325,63563,65463,0),
        (43330,50430,55142,58603,61325,63564,65463,0),
        (43332,50432,55143,58604,61326,63564,65464,0),
        (43334,50433,55144,58605,61326,63565,65464,0),
        (43336,50435,55145,58606,61327,63565,65465,0),
        (43338,50436,55146,58607,61328,63566,65465,0),
        (43340,50438,55147,58607,61328,63566,65466,0),
        (43343,50439,55148,58608,61329,63567,65466,0),
        (43345,50440,55149,58609,61330,63567,65466,0),
        (43347,50441,55150,58609,61330,63568,65467,0),
        (43350,50443,55151,58610,61331,63568,65467,0),
        (43352,50444,55152,58611,61331,63569,65468,0),
        (43353,50445,55153,58612,61332,63569,65468,0),
        (43355,50447,55154,58612,61332,63570,65469,0),
        (43358,50448,55155,58613,61333,63570,65469,0),
        (43360,50450,55156,58614,61334,63571,65469,0),
        (43362,50451,55157,58615,61334,63571,65470,0),
        (43365,50453,55158,58615,61335,63572,65470,0),
        (43367,50454,55159,58616,61335,63572,65471,0),
        (43369,50455,55159,58617,61336,63573,65471,0),
        (43371,50457,55161,58618,61337,63573,65472,0),
        (43373,50458,55162,58618,61337,63574,65472,0),
        (43375,50459,55162,58619,61338,63574,65473,0),
        (43377,50460,55164,58620,61338,63575,65473,0),
        (43380,50462,55165,58620,61339,63575,65473,0),
        (43382,50463,55165,58621,61339,63576,65474,0),
        (43384,50465,55166,58622,61340,63576,65474,0),
        (43386,50466,55168,58623,61341,63577,65475,0),
        (43389,50468,55168,58623,61341,63577,65475,0),
        (43391,50469,55169,58624,61342,63578,65476,0),
        (43393,50470,55170,58625,61343,63578,65476,0),
        (43395,50472,55171,58626,61343,63579,65476,0),
        (43397,50473,55172,58626,61344,63579,65477,0),
        (43399,50474,55173,58627,61344,63580,65477,0),
        (43401,50476,55174,58628,61345,63580,65478,0),
        (43404,50477,55175,58629,61346,63581,65478,0),
        (43406,50478,55176,58629,61346,63581,65479,0),
        (43408,50480,55177,58630,61347,63582,65479,0),
        (43411,50481,55178,58631,61347,63582,65479,0),
        (43413,50483,55179,58631,61348,63583,65480,0),
        (43414,50484,55180,58632,61349,63583,65480,0),
        (43416,50486,55181,58633,61349,63584,65481,0),
        (43419,50487,55182,58634,61350,63584,65481,0),
        (43421,50488,55183,58634,61350,63585,65482,0),
        (43423,50489,55184,58635,61351,63585,65482,0),
        (43426,50491,55185,58636,61352,63586,65482,0),
        (43428,50492,55186,58637,61352,63586,65483,0),
        (43430,50493,55187,58638,61353,63587,65483,0),
        (43432,50495,55188,58638,61353,63587,65484,0),
        (43434,50496,55189,58639,61354,63588,65484,0),
        (43436,50498,55189,58640,61355,63588,65485,0),
        (43438,50499,55191,58641,61355,63589,65485,0),
        (43441,50501,55192,58641,61356,63589,65485,0),
        (43443,50502,55192,58642,61356,63590,65486,0),
        (43445,50503,55193,58643,61357,63590,65486,0),
        (43447,50505,55195,58643,61358,63591,65487,0),
        (43450,50506,55195,58644,61358,63591,65487,0),
        (43451,50507,55196,58645,61359,63592,65488,0),
        (43453,50508,55198,58646,61359,63592,65488,0),
        (43456,50510,55198,58646,61360,63593,65488,0),
        (43458,50511,55199,58647,61360,63593,65489,0),
        (43460,50513,55200,58648,61361,63594,65489,0),
        (43462,50514,55201,58649,61362,63594,65490,0),
        (43465,50516,55202,58649,61362,63595,65490,0),
        (43467,50517,55203,58650,61363,63595,65491,0),
        (43469,50518,55204,58651,61364,63596,65491,0),
        (43471,50520,55205,58652,61364,63596,65491,0),
        (43473,50521,55206,58652,61365,63597,65492,0),
        (43475,50522,55207,58653,61365,63597,65492,0),
        (43477,50524,55208,58654,61366,63598,65493,0),
        (43480,50525,55209,58654,61366,63598,65493,0),
        (43482,50526,55210,58655,61367,63599,65494,0),
        (43484,50527,55211,58656,61368,63599,65494,0),
        (43487,50529,55212,58657,61368,63600,65494,0),
        (43488,50530,55213,58657,61369,63600,65495,0),
        (43490,50532,55214,58658,61370,63601,65495,0),
        (43492,50533,55215,58659,61370,63601,65496,0),
        (43495,50535,55216,58660,61371,63602,65496,0),
        (43497,50536,55216,58660,61371,63602,65497,0),
        (43499,50537,55218,58661,61372,63603,65497,0),
        (43502,50539,55219,58662,61372,63603,65497,0),
        (43504,50540,55219,58663,61373,63604,65498,0),
        (43505,50541,55220,58663,61374,63604,65498,0),
        (43507,50543,55222,58664,61374,63605,65499,0),
        (43510,50544,55222,58665,61375,63605,65499,0),
        (43512,50545,55223,58665,61376,63606,65500,0),
        (43514,50547,55224,58666,61376,63606,65500,0),
        (43517,50548,55225,58667,61377,63607,65500,0),
        (43519,50550,55226,58668,61377,63607,65501,0),
        (43521,50551,55227,58669,61378,63608,65501,0),
        (43522,50553,55228,58669,61378,63608,65502,0),
        (43525,50554,55229,58670,61379,63609,65502,0),
        (43527,50555,55230,58671,61380,63609,65503,0),
        (43529,50556,55231,58672,61380,63610,65503,0),
        (43532,50558,55232,58672,61381,63610,65503,0),
        (43534,50559,55233,58673,61381,63611,65504,0),
        (43536,50560,55234,58674,61382,63611,65504,0),
        (43538,50562,55235,58674,61383,63612,65505,0),
        (43540,50563,55236,58675,61383,63612,65505,0),
        (43542,50564,55237,58676,61384,63613,65506,0),
        (43544,50566,55238,58677,61384,63613,65506,0),
        (43547,50567,55239,58677,61385,63614,65506,0),
        (43549,50569,55240,58678,61385,63614,65507,0),
        (43551,50570,55240,58679,61386,63615,65507,0),
        (43553,50572,55242,58680,61387,63615,65508,0),
        (43556,50573,55243,58680,61387,63616,65508,0),
        (43557,50574,55243,58681,61388,63616,65509,0),
        (43559,50575,55245,58682,61389,63617,65509,0),
        (43562,50577,55246,58682,61389,63617,65509,0),
        (43564,50578,55246,58683,61390,63618,65510,0),
        (43566,50579,55247,58684,61390,63618,65510,0),
        (43568,50581,55248,58685,61391,63619,65511,0),
        (43571,50582,55249,58685,61391,63619,65511,0),
        (43572,50584,55250,58686,61392,63620,65512,0),
        (43574,50585,55251,58687,61393,63620,65512,0),
        (43577,50586,55252,58688,61393,63621,65512,0),
        (43579,50588,55253,58688,61394,63621,65513,0),
        (43581,50589,55254,58689,61395,63622,65513,0),
        (43583,50591,55255,58690,61395,63622,65514,0),
        (43586,50592,55256,58691,61396,63623,65514,0),
        (43588,50593,55257,58691,61396,63623,65515,0),
        (43589,50594,55258,58692,61397,63624,65515,0),
        (43592,50596,55259,58693,61397,63624,65515,0),
        (43594,50597,55260,58693,61398,63625,65516,0),
        (43596,50598,55261,58694,61399,63625,65516,0),
        (43598,50600,55262,58695,61399,63626,65517,0),
        (43601,50601,55263,58696,61400,63626,65517,0),
        (43603,50603,55264,58696,61401,63627,65518,0),
        (43604,50604,55265,58697,61401,63627,65518,0),
        (43607,50606,55266,58698,61402,63628,65518,0),
        (43609,50607,55267,58699,61402,63628,65519,0),
        (43611,50608,55267,58700,61403,63629,65519,0),
        (43613,50610,55269,58700,61403,63629,65520,0),
        (43616,50611,55269,58701,61404,63630,65520,0),
        (43618,50612,55270,58701,61405,63630,65521,0),
        (43620,50613,55272,58702,61405,63631,65521,0),
        (43622,50615,55272,58703,61406,63631,65521,0),
        (43624,50616,55273,58704,61406,63632,65522,0),
        (43626,50617,55274,58705,61407,63632,65522,0),
        (43628,50619,55275,58705,61408,63633,65523,0),
        (43631,50620,55276,58706,61408,63633,65523,0),
        (43633,50622,55277,58707,61409,63634,65524,0),
        (43635,50623,55278,58708,61409,63634,65524,0),
        (43637,50625,55279,58708,61410,63635,65524,0),
        (43639,50626,55280,58709,61410,63635,65525,0),
        (43641,50627,55281,58710,61411,63636,65525,0),
        (43643,50629,55282,58710,61412,63636,65526,0),
        (43646,50630,55283,58711,61412,63637,65526,0),
        (43648,50631,55284,58712,61413,63637,65527,0),
        (43650,50632,55285,58713,61414,63638,65527,0),
        (43652,50634,55286,58713,61414,63638,65527,0),
        (43654,50635,55287,58714,61415,63639,65528,0),
        (43656,50636,55288,58715,61415,63639,65528,0),
        (43658,50638,55289,58716,61416,63640,65529,0),
        (43661,50639,55290,58716,61416,63640,65529,0),
        (43663,50641,55290,58717,61417,63641,65530,0),
        (43665,50642,55292,58718,61418,63641,65530,0),
        (43667,50643,55293,58719,61418,63642,65530,0),
        (43669,50645,55293,58719,61419,63642,65531,0),
        (43671,50646,55294,58720,61419,63643,65531,0),
        (43673,50648,55295,58721,61420,63643,65532,0),
        (43676,50649,55296,58721,61421,63644,65532,0),
        (43678,50650,55297,58722,61421,63644,65533,0),
        (43680,50651,55298,58723,61422,63645,65533,0),
        (43682,50653,55299,58724,61422,63645,65533,0),
        (43684,50654,55300,58724,61423,63646,65534,0),
        (43686,50655,55301,58725,61424,63646,65534,0),
        (43688,50657,55302,58726,61424,63647,65535,0),
        (43690,50658,55303,58726,61424,63647,65535,0)          
);
end TanLROM; 