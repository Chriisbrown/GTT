library ieee;
use ieee.std_logic_1164.all;
use ieee.std_logic_misc.all;
use ieee.numeric_std.all;

package TanLROM is
    type intArray is array(natural range <>) of integer;
    type intArray2D is array(natural range <>) of intArray;


 
     
    constant TanLLUT : intArray(0 to 1023) := (
0,
3,
6,
9,
12,
15,
18,
21,
24,
27,
30,
33,
36,
39,
42,
45,
48,
51,
54,
57,
60,
63,
66,
69,
72,
75,
78,
81,
84,
87,
89,
92,
95,
98,
101,
104,
107,
110,
113,
116,
119,
122,
124,
127,
130,
133,
136,
139,
142,
144,
147,
150,
153,
156,
158,
161,
164,
167,
169,
172,
175,
178,
180,
183,
186,
189,
191,
194,
197,
199,
202,
205,
207,
210,
212,
215,
218,
220,
223,
225,
228,
231,
233,
236,
238,
241,
243,
246,
248,
251,
253,
256,
258,
261,
263,
265,
268,
270,
273,
275,
278,
280,
282,
285,
287,
289,
292,
294,
296,
299,
301,
303,
305,
308,
310,
312,
314,
317,
319,
321,
323,
326,
328,
330,
332,
334,
336,
339,
341,
343,
345,
347,
349,
351,
353,
356,
358,
360,
362,
364,
366,
368,
370,
372,
374,
376,
378,
380,
382,
384,
386,
388,
390,
392,
394,
396,
397,
399,
401,
403,
405,
407,
409,
411,
413,
414,
416,
418,
420,
422,
424,
425,
427,
429,
431,
433,
434,
436,
438,
440,
441,
443,
445,
447,
448,
450,
452,
454,
455,
457,
459,
460,
462,
464,
465,
467,
469,
470,
472,
474,
475,
477,
479,
480,
482,
483,
485,
487,
488,
490,
491,
493,
494,
496,
498,
499,
501,
502,
504,
505,
507,
508,
510,
511,
513,
514,
516,
517,
519,
520,
522,
523,
525,
526,
528,
529,
530,
532,
533,
535,
536,
538,
539,
540,
542,
543,
545,
546,
547,
549,
550,
552,
553,
554,
556,
557,
558,
560,
561,
562,
564,
565,
566,
568,
569,
570,
572,
573,
574,
576,
577,
578,
579,
581,
582,
583,
585,
586,
587,
588,
590,
591,
592,
593,
595,
596,
597,
598,
600,
601,
602,
603,
604,
606,
607,
608,
609,
611,
612,
613,
614,
615,
616,
618,
619,
620,
621,
622,
623,
625,
626,
627,
628,
629,
630,
632,
633,
634,
635,
636,
637,
638,
639,
641,
642,
643,
644,
645,
646,
647,
648,
649,
650,
652,
653,
654,
655,
656,
657,
658,
659,
660,
661,
662,
663,
664,
665,
666,
667,
669,
670,
671,
672,
673,
674,
675,
676,
677,
678,
679,
680,
681,
682,
683,
684,
685,
686,
687,
688,
689,
690,
691,
692,
693,
694,
695,
696,
697,
698,
699,
700,
701,
701,
702,
703,
704,
705,
706,
707,
708,
709,
710,
711,
712,
713,
714,
715,
716,
717,
718,
718,
719,
720,
721,
722,
723,
724,
725,
726,
727,
728,
728,
729,
730,
731,
732,
733,
734,
735,
736,
736,
737,
738,
739,
740,
741,
742,
743,
743,
744,
745,
746,
747,
748,
749,
749,
750,
751,
752,
753,
754,
755,
755,
756,
757,
758,
759,
760,
760,
761,
762,
763,
764,
765,
765,
766,
767,
768,
769,
769,
770,
771,
772,
773,
773,
774,
775,
776,
777,
777,
778,
779,
780,
781,
781,
782,
783,
784,
785,
785,
786,
787,
788,
788,
789,
790,
791,
792,
792,
793,
794,
795,
795,
796,
797,
798,
798,
799,
800,
801,
801,
802,
803,
804,
804,
805,
806,
807,
807,
808,
809,
810,
810,
811,
812,
812,
813,
814,
815,
815,
816,
817,
818,
818,
819,
820,
820,
821,
822,
823,
823,
824,
825,
825,
826,
827,
828,
828,
829,
830,
830,
831,
832,
832,
833,
834,
834,
835,
836,
837,
837,
838,
839,
839,
840,
841,
841,
842,
843,
843,
844,
845,
845,
846,
847,
847,
848,
849,
849,
850,
851,
851,
852,
853,
853,
854,
855,
855,
856,
857,
857,
858,
859,
859,
860,
861,
861,
862,
862,
863,
864,
864,
865,
866,
866,
867,
868,
868,
869,
869,
870,
871,
871,
872,
873,
873,
874,
874,
875,
876,
876,
877,
878,
878,
879,
879,
880,
881,
881,
882,
883,
883,
884,
884,
885,
886,
886,
887,
887,
888,
889,
889,
890,
890,
891,
892,
892,
893,
893,
894,
895,
895,
896,
896,
897,
897,
898,
899,
899,
900,
900,
901,
902,
902,
903,
903,
904,
904,
905,
906,
906,
907,
907,
908,
909,
909,
910,
910,
911,
911,
912,
913,
913,
914,
914,
915,
915,
916,
916,
917,
918,
918,
919,
919,
920,
920,
921,
921,
922,
923,
923,
924,
924,
925,
925,
926,
926,
927,
928,
928,
929,
929,
930,
930,
931,
931,
932,
932,
933,
933,
934,
935,
935,
936,
936,
937,
937,
938,
938,
939,
939,
940,
940,
941,
941,
942,
942,
943,
944,
944,
945,
945,
946,
946,
947,
947,
948,
948,
949,
949,
950,
950,
951,
951,
952,
952,
953,
953,
954,
954,
955,
955,
956,
956,
957,
957,
958,
958,
959,
959,
960,
960,
961,
961,
962,
962,
963,
963,
964,
964,
965,
965,
966,
966,
967,
967,
968,
968,
969,
969,
970,
970,
971,
971,
972,
972,
973,
973,
974,
974,
975,
975,
976,
976,
977,
977,
978,
978,
979,
979,
980,
980,
980,
981,
981,
982,
982,
983,
983,
984,
984,
985,
985,
986,
986,
987,
987,
988,
988,
988,
989,
989,
990,
990,
991,
991,
992,
992,
993,
993,
994,
994,
995,
995,
995,
996,
996,
997,
997,
998,
998,
999,
999,
1000,
1000,
1000,
1001,
1001,
1002,
1002,
1003,
1003,
1004,
1004,
1004,
1005,
1005,
1006,
1006,
1007,
1007,
1008,
1008,
1009,
1009,
1009,
1010,
1010,
1011,
1011,
1012,
1012,
1012,
1013,
1013,
1014,
1014,
1015,
1015,
1016,
1016,
1016,
1017,
1017,
1018,
1018,
1019,
1019,
1019,
1020,
1020,
1021,
1021,
1022,
1022,
1022,
1023,
1023,
1024,
1024,
1025,
1025,
1025,
1026,
1026,
1027,
1027,
1028,
1028,
1028,
1029,
1029,
1030,
1030,
1030,
1031,
1031,
1032,
1032,
1033,
1033,
1033,
1034,
1034,
1035,
1035,
1035,
1036,
1036,
1037,
1037,
1038,
1038,
1038,
1039,
1039,
1040,
1040,
1040,
1041,
1041,
1042,
1042,
1042,
1043,
1043,
1044,
1044,
1044,
1045,
1045,
1046,
1046,
1047,
1047,
1047,
1048,
1048,
1049,
1049,
1049,
1050,
1050,
1051,
1051,
1051,
1052,
1052,
1052,
1053,
1053,
1054,
1054,
1054,
1055,
1055,
1056,
1056,
1056,
1057,
1057,
1058,
1058,
1058,
1059,
1059,
1060,
1060,
1060,
1061,
1061,
1062,
1062,
1062,
1063,
1063,
1063,
1064,
1064,
1065,
1065,
1065,
1066,
1066,
1067,
1067,
1067,
1068,
1068,
1068,
1069,
1069,
1070,
1070,
1070,
1071,
1071,
1071,
1072,
1072,
1073,
1073,
1073,
1074        
);


end TanLROM; 