library ieee;
use ieee.std_logic_1164.all;
use ieee.std_logic_misc.all;
use ieee.numeric_std.all;


package ROMConstants is
  type intArray is array(natural range <>) of integer;

  constant TrigArray : intArray(0 TO 194) := (
  255,
  255,
  255,
  255,
  255,
  255,
  255,
  255,
  254,
  254,
  254,
  254,
  254,
  254,
  253,
  253,
  253,
  253,
  252,
  252,
  252,
  251,
  251,
  251,
  250,
  250,
  249,
  249,
  248,
  248,
  248,
  247,
  246,
  246,
  245,
  245,
  244,
  244,
  243,
  242,
  242,
  241,
  240,
  240,
  239,
  238,
  238,
  237,
  236,
  235,
  234,
  234,
  233,
  232,
  231,
  230,
  229,
  228,
  227,
  226,
  225,
  225,
  224,
  223,
  222,
  220,
  219,
  218,
  217,
  216,
  215,
  214,
  213,
  212,
  211,
  209,
  208,
  207,
  206,
  205,
  203,
  202,
  201,
  200,
  198,
  197,
  196,
  194,
  193,
  192,
  190,
  189,
  187,
  186,
  185,
  183,
  182,
  180,
  179,
  177,
  176,
  174,
  173,
  171,
  170,
  168,
  167,
  165,
  164,
  162,
  160,
  159,
  157,
  156,
  154,
  152,
  151,
  149,
  147,
  146,
  144,
  142,
  140,
  139,
  137,
  135,
  133,
  132,
  130,
  128,
  126,
  125,
  123,
  121,
  119,
  117,
  115,
  114,
  112,
  110,
  108,
  106,
  104,
  102,
  100,
  99,
  97,
  95,
  93,
  91,
  89,
  87,
  85,
  83,
  81,
  79,
  77,
  75,
  73,
  71,
  69,
  67,
  65,
  63,
  61,
  59,
  57,
  55,
  53,
  51,
  49,
  47,
  45,
  43,
  41,
  39,
  37,
  35,
  33,
  31,
  29,
  27,
  25,
  23,
  21,
  19,
  17,
  14,
  12,
  10,
  8,
  6,
  4,
  2,
  0);


end ROMConstants;
  